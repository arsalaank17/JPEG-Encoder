-- Automatically generated VHDL-93
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;
use std.textio.all;
use work.all;
use work.Main_topEntity_types.all;

entity topEntity is
  port(input_0_0 : in signed(63 downto 0);
       input_0_1 : in signed(63 downto 0);
       input_0_2 : in signed(63 downto 0);
       input_0_3 : in signed(63 downto 0);
       input_0_4 : in signed(63 downto 0);
       input_0_5 : in signed(63 downto 0);
       input_0_6 : in signed(63 downto 0);
       input_0_7 : in signed(63 downto 0);
       input_1_0 : in signed(63 downto 0);
       input_1_1 : in signed(63 downto 0);
       input_1_2 : in signed(63 downto 0);
       input_1_3 : in signed(63 downto 0);
       input_1_4 : in signed(63 downto 0);
       input_1_5 : in signed(63 downto 0);
       input_1_6 : in signed(63 downto 0);
       input_1_7 : in signed(63 downto 0);
       input_2_0 : in signed(63 downto 0);
       input_2_1 : in signed(63 downto 0);
       input_2_2 : in signed(63 downto 0);
       input_2_3 : in signed(63 downto 0);
       input_2_4 : in signed(63 downto 0);
       input_2_5 : in signed(63 downto 0);
       input_2_6 : in signed(63 downto 0);
       input_2_7 : in signed(63 downto 0);
       input_3_0 : in signed(63 downto 0);
       input_3_1 : in signed(63 downto 0);
       input_3_2 : in signed(63 downto 0);
       input_3_3 : in signed(63 downto 0);
       input_3_4 : in signed(63 downto 0);
       input_3_5 : in signed(63 downto 0);
       input_3_6 : in signed(63 downto 0);
       input_3_7 : in signed(63 downto 0);
       input_4_0 : in signed(63 downto 0);
       input_4_1 : in signed(63 downto 0);
       input_4_2 : in signed(63 downto 0);
       input_4_3 : in signed(63 downto 0);
       input_4_4 : in signed(63 downto 0);
       input_4_5 : in signed(63 downto 0);
       input_4_6 : in signed(63 downto 0);
       input_4_7 : in signed(63 downto 0);
       input_5_0 : in signed(63 downto 0);
       input_5_1 : in signed(63 downto 0);
       input_5_2 : in signed(63 downto 0);
       input_5_3 : in signed(63 downto 0);
       input_5_4 : in signed(63 downto 0);
       input_5_5 : in signed(63 downto 0);
       input_5_6 : in signed(63 downto 0);
       input_5_7 : in signed(63 downto 0);
       input_6_0 : in signed(63 downto 0);
       input_6_1 : in signed(63 downto 0);
       input_6_2 : in signed(63 downto 0);
       input_6_3 : in signed(63 downto 0);
       input_6_4 : in signed(63 downto 0);
       input_6_5 : in signed(63 downto 0);
       input_6_6 : in signed(63 downto 0);
       input_6_7 : in signed(63 downto 0);
       input_7_0 : in signed(63 downto 0);
       input_7_1 : in signed(63 downto 0);
       input_7_2 : in signed(63 downto 0);
       input_7_3 : in signed(63 downto 0);
       input_7_4 : in signed(63 downto 0);
       input_7_5 : in signed(63 downto 0);
       input_7_6 : in signed(63 downto 0);
       input_7_7 : in signed(63 downto 0);
       result_0  : out Main_topEntity_types.Maybe;
       result_1  : out Main_topEntity_types.Maybe;
       result_2  : out Main_topEntity_types.Maybe;
       result_3  : out Main_topEntity_types.Maybe;
       result_4  : out Main_topEntity_types.Maybe;
       result_5  : out Main_topEntity_types.Maybe;
       result_6  : out Main_topEntity_types.Maybe;
       result_7  : out Main_topEntity_types.Maybe;
       result_8  : out Main_topEntity_types.Maybe;
       result_9  : out Main_topEntity_types.Maybe;
       result_10 : out Main_topEntity_types.Maybe;
       result_11 : out Main_topEntity_types.Maybe;
       result_12 : out Main_topEntity_types.Maybe;
       result_13 : out Main_topEntity_types.Maybe;
       result_14 : out Main_topEntity_types.Maybe;
       result_15 : out Main_topEntity_types.Maybe;
       result_16 : out Main_topEntity_types.Maybe;
       result_17 : out Main_topEntity_types.Maybe;
       result_18 : out Main_topEntity_types.Maybe;
       result_19 : out Main_topEntity_types.Maybe;
       result_20 : out Main_topEntity_types.Maybe;
       result_21 : out Main_topEntity_types.Maybe;
       result_22 : out Main_topEntity_types.Maybe;
       result_23 : out Main_topEntity_types.Maybe;
       result_24 : out Main_topEntity_types.Maybe;
       result_25 : out Main_topEntity_types.Maybe;
       result_26 : out Main_topEntity_types.Maybe;
       result_27 : out Main_topEntity_types.Maybe;
       result_28 : out Main_topEntity_types.Maybe;
       result_29 : out Main_topEntity_types.Maybe;
       result_30 : out Main_topEntity_types.Maybe;
       result_31 : out Main_topEntity_types.Maybe;
       result_32 : out Main_topEntity_types.Maybe;
       result_33 : out Main_topEntity_types.Maybe;
       result_34 : out Main_topEntity_types.Maybe;
       result_35 : out Main_topEntity_types.Maybe;
       result_36 : out Main_topEntity_types.Maybe;
       result_37 : out Main_topEntity_types.Maybe;
       result_38 : out Main_topEntity_types.Maybe;
       result_39 : out Main_topEntity_types.Maybe;
       result_40 : out Main_topEntity_types.Maybe;
       result_41 : out Main_topEntity_types.Maybe;
       result_42 : out Main_topEntity_types.Maybe;
       result_43 : out Main_topEntity_types.Maybe;
       result_44 : out Main_topEntity_types.Maybe;
       result_45 : out Main_topEntity_types.Maybe;
       result_46 : out Main_topEntity_types.Maybe;
       result_47 : out Main_topEntity_types.Maybe;
       result_48 : out Main_topEntity_types.Maybe;
       result_49 : out Main_topEntity_types.Maybe;
       result_50 : out Main_topEntity_types.Maybe;
       result_51 : out Main_topEntity_types.Maybe;
       result_52 : out Main_topEntity_types.Maybe;
       result_53 : out Main_topEntity_types.Maybe;
       result_54 : out Main_topEntity_types.Maybe;
       result_55 : out Main_topEntity_types.Maybe;
       result_56 : out Main_topEntity_types.Maybe;
       result_57 : out Main_topEntity_types.Maybe;
       result_58 : out Main_topEntity_types.Maybe;
       result_59 : out Main_topEntity_types.Maybe;
       result_60 : out Main_topEntity_types.Maybe;
       result_61 : out Main_topEntity_types.Maybe;
       result_62 : out Main_topEntity_types.Maybe;
       result_63 : out Main_topEntity_types.Maybe);
end;

architecture structural of topEntity is
  signal \c$app_arg\                : Main_topEntity_types.array_of_signed_64(0 to 63);
  signal result_128                 : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out\                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg\         : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2                         : signed(63 downto 0);
  signal \c$~<~Out_app_arg_0\       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_0                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y                          : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_1                       : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut\      : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes                    : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr                     : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_0\    : boolean;
  signal \c$~<~Out_app_arg_1\       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_0                        : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1                         : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2                      : signed(63 downto 0);
  signal \c$countConOut_app_arg\    : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_0\               : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_2\       : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_2                       : signed(63 downto 0);
  signal \c$~<~Out_case_alt\        : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_3                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_1                        : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1                         : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_1\    : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_0                  : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_0                   : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_2\    : boolean;
  signal \c$~<~Out_app_arg_3\       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_2                        : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_0                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_0                    : signed(63 downto 0);
  signal \c$countConOut_app_arg_0\  : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_1\               : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_4\       : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_4                       : signed(63 downto 0);
  signal \c$~<~Out_case_alt_0\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_5                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_3                        : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_0                       : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_3\    : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_1                  : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_1                   : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_4\    : boolean;
  signal \c$~<~Out_app_arg_5\       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_4                        : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_1                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_1                    : signed(63 downto 0);
  signal \c$countConOut_app_arg_1\  : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_2\               : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_6\       : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_6                       : signed(63 downto 0);
  signal \c$~<~Out_case_alt_1\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_7                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_5                        : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_1                       : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_5\    : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_2                  : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_2                   : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_6\    : boolean;
  signal \c$~<~Out_app_arg_7\       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_6                        : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_2                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_2                    : signed(63 downto 0);
  signal \c$countConOut_app_arg_2\  : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_3\               : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_8\       : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_8                       : signed(63 downto 0);
  signal \c$~<~Out_case_alt_2\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_9                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_7                        : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_2                       : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_7\    : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_3                  : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_3                   : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_8\    : boolean;
  signal \c$~<~Out_app_arg_9\       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_8                        : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_3                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_3                    : signed(63 downto 0);
  signal \c$countConOut_app_arg_3\  : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_4\               : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_10\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_10                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_3\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_11                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_9                        : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_3                       : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_9\    : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_4                  : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_4                   : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_10\   : boolean;
  signal \c$~<~Out_app_arg_11\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_10                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_4                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_4                    : signed(63 downto 0);
  signal \c$countConOut_app_arg_4\  : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_5\               : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_12\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_12                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_4\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_13                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_11                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_4                       : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_11\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_5                  : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_5                   : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_12\   : boolean;
  signal \c$~<~Out_app_arg_13\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_12                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_5                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_5                    : signed(63 downto 0);
  signal \c$countConOut_app_arg_5\  : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_6\               : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_14\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_14                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_5\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_15                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_13                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_5                       : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_13\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_6                  : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_6                   : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_14\   : boolean;
  signal \c$~<~Out_app_arg_15\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_14                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_6                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_6                    : signed(63 downto 0);
  signal \c$countConOut_app_arg_6\  : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_7\               : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_16\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_16                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_6\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_17                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_15                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_6                       : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_15\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_7                  : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_7                   : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_16\   : boolean;
  signal \c$~<~Out_app_arg_17\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_16                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_7                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_7                    : signed(63 downto 0);
  signal \c$countConOut_app_arg_7\  : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_8\               : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_18\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_18                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_7\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_19                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_17                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_7                       : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_17\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_8                  : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_8                   : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_18\   : boolean;
  signal \c$~<~Out_app_arg_19\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_18                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_8                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_8                    : signed(63 downto 0);
  signal \c$countConOut_app_arg_8\  : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_9\               : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_20\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_20                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_8\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_21                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_19                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_8                       : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_19\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_9                  : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_9                   : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_20\   : boolean;
  signal \c$~<~Out_app_arg_21\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_20                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_9                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_9                    : signed(63 downto 0);
  signal \c$countConOut_app_arg_9\  : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_10\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_22\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_22                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_9\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_23                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_21                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_9                       : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_21\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_10                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_10                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_22\   : boolean;
  signal \c$~<~Out_app_arg_23\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_22                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_10                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_10                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_10\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_11\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_24\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_24                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_10\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_25                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_23                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_10                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_23\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_11                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_11                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_24\   : boolean;
  signal \c$~<~Out_app_arg_25\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_24                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_11                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_11                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_11\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_12\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_26\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_26                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_11\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_27                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_25                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_11                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_25\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_12                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_12                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_26\   : boolean;
  signal \c$~<~Out_app_arg_27\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_26                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_12                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_12                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_12\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_13\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_28\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_28                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_12\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_29                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_27                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_12                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_27\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_13                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_13                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_28\   : boolean;
  signal \c$~<~Out_app_arg_29\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_28                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_13                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_13                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_13\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_14\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_30\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_30                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_13\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_31                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_29                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_13                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_29\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_14                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_14                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_30\   : boolean;
  signal \c$~<~Out_app_arg_31\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_30                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_14                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_14                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_14\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_15\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_32\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_32                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_14\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_33                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_31                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_14                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_31\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_15                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_15                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_32\   : boolean;
  signal \c$~<~Out_app_arg_33\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_32                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_15                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_15                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_15\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_16\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_34\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_34                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_15\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_35                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_33                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_15                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_33\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_16                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_16                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_34\   : boolean;
  signal \c$~<~Out_app_arg_35\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_34                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_16                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_16                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_16\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_17\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_36\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_36                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_16\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_37                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_35                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_16                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_35\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_17                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_17                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_36\   : boolean;
  signal \c$~<~Out_app_arg_37\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_36                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_17                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_17                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_17\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_18\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_38\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_38                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_17\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_39                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_37                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_17                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_37\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_18                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_18                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_38\   : boolean;
  signal \c$~<~Out_app_arg_39\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_38                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_18                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_18                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_18\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_19\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_40\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_40                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_18\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_41                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_39                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_18                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_39\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_19                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_19                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_40\   : boolean;
  signal \c$~<~Out_app_arg_41\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_40                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_19                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_19                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_19\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_20\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_42\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_42                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_19\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_43                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_41                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_19                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_41\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_20                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_20                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_42\   : boolean;
  signal \c$~<~Out_app_arg_43\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_42                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_20                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_20                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_20\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_21\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_44\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_44                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_20\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_45                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_43                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_20                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_43\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_21                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_21                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_44\   : boolean;
  signal \c$~<~Out_app_arg_45\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_44                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_21                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_21                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_21\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_22\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_46\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_46                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_21\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_47                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_45                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_21                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_45\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_22                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_22                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_46\   : boolean;
  signal \c$~<~Out_app_arg_47\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_46                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_22                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_22                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_22\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_23\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_48\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_48                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_22\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_49                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_47                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_22                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_47\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_23                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_23                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_48\   : boolean;
  signal \c$~<~Out_app_arg_49\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_48                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_23                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_23                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_23\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_24\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_50\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_50                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_23\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_51                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_49                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_23                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_49\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_24                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_24                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_50\   : boolean;
  signal \c$~<~Out_app_arg_51\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_50                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_24                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_24                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_24\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_25\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_52\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_52                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_24\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_53                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_51                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_24                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_51\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_25                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_25                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_52\   : boolean;
  signal \c$~<~Out_app_arg_53\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_52                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_25                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_25                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_25\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_26\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_54\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_54                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_25\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_55                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_53                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_25                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_53\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_26                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_26                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_54\   : boolean;
  signal \c$~<~Out_app_arg_55\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_54                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_26                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_26                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_26\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_27\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_56\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_56                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_26\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_57                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_55                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_26                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_55\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_27                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_27                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_56\   : boolean;
  signal \c$~<~Out_app_arg_57\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_56                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_27                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_27                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_27\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_28\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_58\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_58                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_27\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_59                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_57                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_27                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_57\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_28                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_28                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_58\   : boolean;
  signal \c$~<~Out_app_arg_59\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_58                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_28                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_28                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_28\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_29\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_60\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_60                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_28\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_61                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_59                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_28                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_59\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_29                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_29                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_60\   : boolean;
  signal \c$~<~Out_app_arg_61\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_60                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_29                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_29                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_29\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_30\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_62\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_62                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_29\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_63                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_61                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_29                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_61\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_30                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_30                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_62\   : boolean;
  signal \c$~<~Out_app_arg_63\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_62                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_30                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_30                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_30\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_31\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_64\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_64                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_30\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_65                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_63                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_30                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_63\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_31                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_31                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_64\   : boolean;
  signal \c$~<~Out_app_arg_65\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_64                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_31                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_31                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_31\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_32\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_66\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_66                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_31\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_67                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_65                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_31                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_65\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_32                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_32                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_66\   : boolean;
  signal \c$~<~Out_app_arg_67\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_66                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_32                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_32                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_32\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_33\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_68\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_68                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_32\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_69                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_67                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_32                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_67\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_33                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_33                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_68\   : boolean;
  signal \c$~<~Out_app_arg_69\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_68                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_33                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_33                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_33\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_34\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_70\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_70                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_33\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_71                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_69                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_33                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_69\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_34                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_34                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_70\   : boolean;
  signal \c$~<~Out_app_arg_71\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_70                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_34                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_34                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_34\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_35\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_72\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_72                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_34\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_73                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_71                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_34                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_71\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_35                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_35                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_72\   : boolean;
  signal \c$~<~Out_app_arg_73\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_72                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_35                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_35                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_35\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_36\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_74\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_74                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_35\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_75                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_73                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_35                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_73\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_36                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_36                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_74\   : boolean;
  signal \c$~<~Out_app_arg_75\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_74                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_36                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_36                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_36\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_37\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_76\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_76                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_36\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_77                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_75                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_36                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_75\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_37                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_37                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_76\   : boolean;
  signal \c$~<~Out_app_arg_77\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_76                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_37                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_37                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_37\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_38\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_78\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_78                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_37\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_79                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_77                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_37                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_77\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_38                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_38                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_78\   : boolean;
  signal \c$~<~Out_app_arg_79\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_78                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_38                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_38                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_38\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_39\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_80\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_80                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_38\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_81                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_79                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_38                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_79\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_39                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_39                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_80\   : boolean;
  signal \c$~<~Out_app_arg_81\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_80                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_39                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_39                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_39\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_40\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_82\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_82                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_39\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_83                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_81                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_39                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_81\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_40                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_40                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_82\   : boolean;
  signal \c$~<~Out_app_arg_83\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_82                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_40                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_40                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_40\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_41\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_84\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_84                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_40\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_85                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_83                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_40                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_83\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_41                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_41                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_84\   : boolean;
  signal \c$~<~Out_app_arg_85\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_84                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_41                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_41                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_41\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_42\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_86\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_86                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_41\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_87                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_85                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_41                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_85\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_42                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_42                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_86\   : boolean;
  signal \c$~<~Out_app_arg_87\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_86                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_42                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_42                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_42\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_43\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_88\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_88                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_42\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_89                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_87                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_42                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_87\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_43                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_43                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_88\   : boolean;
  signal \c$~<~Out_app_arg_89\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_88                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_43                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_43                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_43\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_44\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_90\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_90                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_43\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_91                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_89                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_43                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_89\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_44                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_44                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_90\   : boolean;
  signal \c$~<~Out_app_arg_91\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_90                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_44                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_44                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_44\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_45\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_92\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_92                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_44\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_93                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_91                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_44                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_91\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_45                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_45                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_92\   : boolean;
  signal \c$~<~Out_app_arg_93\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_92                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_45                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_45                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_45\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_46\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_94\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_94                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_45\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_95                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_93                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_45                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_93\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_46                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_46                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_94\   : boolean;
  signal \c$~<~Out_app_arg_95\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_94                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_46                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_46                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_46\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_47\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_96\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_96                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_46\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_97                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_95                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_46                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_95\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_47                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_47                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_96\   : boolean;
  signal \c$~<~Out_app_arg_97\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_96                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_47                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_47                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_47\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_48\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_98\      : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_98                      : signed(63 downto 0);
  signal \c$~<~Out_case_alt_47\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_99                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_97                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_47                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_97\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_48                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_48                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_98\   : boolean;
  signal \c$~<~Out_app_arg_99\      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_98                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_48                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_48                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_48\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_49\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_100\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_100                     : signed(63 downto 0);
  signal \c$~<~Out_case_alt_48\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_101                     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_99                       : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_48                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_99\   : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_49                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_49                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_100\  : boolean;
  signal \c$~<~Out_app_arg_101\     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_100                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_49                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_49                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_49\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_50\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_102\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_102                     : signed(63 downto 0);
  signal \c$~<~Out_case_alt_49\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_103                     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_101                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_49                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_101\  : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_50                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_50                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_102\  : boolean;
  signal \c$~<~Out_app_arg_103\     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_102                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_50                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_50                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_50\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_51\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_104\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_104                     : signed(63 downto 0);
  signal \c$~<~Out_case_alt_50\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_105                     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_103                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_50                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_103\  : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_51                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_51                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_104\  : boolean;
  signal \c$~<~Out_app_arg_105\     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_104                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_51                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_51                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_51\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_52\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_106\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_106                     : signed(63 downto 0);
  signal \c$~<~Out_case_alt_51\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_107                     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_105                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_51                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_105\  : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_52                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_52                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_106\  : boolean;
  signal \c$~<~Out_app_arg_107\     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_106                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_52                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_52                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_52\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_53\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_108\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_108                     : signed(63 downto 0);
  signal \c$~<~Out_case_alt_52\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_109                     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_107                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_52                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_107\  : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_53                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_53                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_108\  : boolean;
  signal \c$~<~Out_app_arg_109\     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_108                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_53                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_53                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_53\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_54\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_110\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_110                     : signed(63 downto 0);
  signal \c$~<~Out_case_alt_53\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_111                     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_109                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_53                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_109\  : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_54                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_54                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_110\  : boolean;
  signal \c$~<~Out_app_arg_111\     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_110                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_54                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_54                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_54\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_55\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_112\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_112                     : signed(63 downto 0);
  signal \c$~<~Out_case_alt_54\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_113                     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_111                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_54                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_111\  : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_55                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_55                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_112\  : boolean;
  signal \c$~<~Out_app_arg_113\     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_112                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_55                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_55                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_55\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_56\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_114\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_114                     : signed(63 downto 0);
  signal \c$~<~Out_case_alt_55\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_115                     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_113                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_55                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_113\  : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_56                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_56                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_114\  : boolean;
  signal \c$~<~Out_app_arg_115\     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_114                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_56                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_56                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_56\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_57\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_116\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_116                     : signed(63 downto 0);
  signal \c$~<~Out_case_alt_56\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_117                     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_115                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_56                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_115\  : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_57                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_57                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_116\  : boolean;
  signal \c$~<~Out_app_arg_117\     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_116                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_57                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_57                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_57\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_58\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_118\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_118                     : signed(63 downto 0);
  signal \c$~<~Out_case_alt_57\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_119                     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_117                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_57                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_117\  : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_58                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_58                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_118\  : boolean;
  signal \c$~<~Out_app_arg_119\     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_118                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_58                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_58                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_58\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_59\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_120\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_120                     : signed(63 downto 0);
  signal \c$~<~Out_case_alt_58\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_121                     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_119                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_58                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_119\  : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_59                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_59                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_120\  : boolean;
  signal \c$~<~Out_app_arg_121\     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_120                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_59                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_59                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_59\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_60\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_122\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_122                     : signed(63 downto 0);
  signal \c$~<~Out_case_alt_59\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_123                     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_121                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_59                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_121\  : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_60                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_60                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_122\  : boolean;
  signal \c$~<~Out_app_arg_123\     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_122                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_60                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_60                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_60\ : Main_topEntity_types.Tup2_0;
  signal \c$~<~Out_61\              : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$~<~Out_app_arg_124\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_124                     : signed(63 downto 0);
  signal \c$~<~Out_case_alt_60\     : Main_topEntity_types.Tup2;
  -- Run-Length-Encoding.hs:50:1-8
  signal x2_125                     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_123                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal a1_60                      : Main_topEntity_types.Tup2_1;
  signal \c$~<~Out_case_scrut_123\  : Main_topEntity_types.Maybe;
  -- Run-Length-Encoding.hs:50:1-8
  signal currRes_61                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  -- Run-Length-Encoding.hs:50:1-8
  signal resPtr_61                  : signed(63 downto 0);
  signal \c$~<~Out_case_scrut_124\  : boolean;
  signal \c$~<~Out_app_arg_125\     : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal y_124                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_61                      : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_61                   : signed(63 downto 0);
  signal \c$countConOut_app_arg_61\ : signed(63 downto 0);
  signal result_129                 : Main_topEntity_types.array_of_Maybe(0 to 63);
  signal \c$countConOut_case_scrut\ : boolean;
  signal \c$countConOut_app_arg_62\ : Main_topEntity_types.Tup2_0;
  -- Run-Length-Encoding.hs:50:1-8
  signal wild2_62                   : signed(63 downto 0);
  -- Run-Length-Encoding.hs:50:1-8
  signal x1_62                      : signed(63 downto 0);
  signal r_input                    : Main_topEntity_types.array_of_array_of_8_signed_64(0 to 7);
  signal result                     : Main_topEntity_types.array_of_Maybe(0 to 63);

begin
  r_input <= Main_topEntity_types.array_of_array_of_8_signed_64'( Main_topEntity_types.array_of_signed_64'( input_0_0
                                                                                                          , input_0_1
                                                                                                          , input_0_2
                                                                                                          , input_0_3
                                                                                                          , input_0_4
                                                                                                          , input_0_5
                                                                                                          , input_0_6
                                                                                                          , input_0_7 )
                                                                , Main_topEntity_types.array_of_signed_64'( input_1_0
                                                                                                          , input_1_1
                                                                                                          , input_1_2
                                                                                                          , input_1_3
                                                                                                          , input_1_4
                                                                                                          , input_1_5
                                                                                                          , input_1_6
                                                                                                          , input_1_7 )
                                                                , Main_topEntity_types.array_of_signed_64'( input_2_0
                                                                                                          , input_2_1
                                                                                                          , input_2_2
                                                                                                          , input_2_3
                                                                                                          , input_2_4
                                                                                                          , input_2_5
                                                                                                          , input_2_6
                                                                                                          , input_2_7 )
                                                                , Main_topEntity_types.array_of_signed_64'( input_3_0
                                                                                                          , input_3_1
                                                                                                          , input_3_2
                                                                                                          , input_3_3
                                                                                                          , input_3_4
                                                                                                          , input_3_5
                                                                                                          , input_3_6
                                                                                                          , input_3_7 )
                                                                , Main_topEntity_types.array_of_signed_64'( input_4_0
                                                                                                          , input_4_1
                                                                                                          , input_4_2
                                                                                                          , input_4_3
                                                                                                          , input_4_4
                                                                                                          , input_4_5
                                                                                                          , input_4_6
                                                                                                          , input_4_7 )
                                                                , Main_topEntity_types.array_of_signed_64'( input_5_0
                                                                                                          , input_5_1
                                                                                                          , input_5_2
                                                                                                          , input_5_3
                                                                                                          , input_5_4
                                                                                                          , input_5_5
                                                                                                          , input_5_6
                                                                                                          , input_5_7 )
                                                                , Main_topEntity_types.array_of_signed_64'( input_6_0
                                                                                                          , input_6_1
                                                                                                          , input_6_2
                                                                                                          , input_6_3
                                                                                                          , input_6_4
                                                                                                          , input_6_5
                                                                                                          , input_6_6
                                                                                                          , input_6_7 )
                                                                , Main_topEntity_types.array_of_signed_64'( input_7_0
                                                                                                          , input_7_1
                                                                                                          , input_7_2
                                                                                                          , input_7_3
                                                                                                          , input_7_4
                                                                                                          , input_7_5
                                                                                                          , input_7_6
                                                                                                          , input_7_7 ) );

  matrixTraversalZigZag1_capp_arg : entity matrixTraversalZigZag1
    port map
      (result  => \c$app_arg\, \input\ => r_input);

  result_128 <= ( Tup2_0_sel0_signed => x2 + to_signed(1,64)
                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out\ ) when \c$~<~Out_case_scrut_0\ else
                ( Tup2_0_sel0_signed => resPtr
                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out\ );

  clash_internal_cOut : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out\
      , xs           => currRes
      , ds           => \c$~<~Out_app_arg\ );

  \c$~<~Out_app_arg\ <= ( Tup2_sel0_signed => x2 + to_signed(1,64)
                        , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2)
                         & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_0\ else
                        ( Tup2_sel0_signed => resPtr
                        , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_0)
                         & std_logic_vector(\c$~<~Out_app_arg_0\)))) );

  x2 <= resPtr;

  with (\c$~<~Out_case_scrut\(128 downto 128)) select
    \c$~<~Out_app_arg_0\ <= signed'(0 to 63 => '-') when "0",
                            x2_0 + to_signed(1,64) when others;

  x2_0 <= y;

  y <= x2_1.Tup2_1_sel1_signed_1;

  x2_1 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut\(127 downto 0)));

  -- index begin
  indexVec : block
    signal vec_index : integer range 0 to 64-1;
  begin
    vec_index <= to_integer(resPtr)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut\ <= currRes(vec_index);
  end block;
  -- index end

  currRes <= \c$countConOut_app_arg\.Tup2_0_sel1_array_of_Maybe;

  resPtr <= \c$countConOut_app_arg\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_0\ <= tagToEnum(\c$~<~Out_app_arg_1\);

  \c$~<~Out_app_arg_1\ <= to_signed(1,64) when x1 /= y_0 else to_signed(0,64);

  y_0 <= wild2_0;

  x1 <= wild2;

  -- index begin
  indexVec_0 : block
    signal vec_index_0 : integer range 0 to 64-1;
  begin
    vec_index_0 <= to_integer(to_signed(63,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2 <= \c$app_arg\(vec_index_0);
  end block;
  -- index end

  \c$countConOut_app_arg\ <= ( Tup2_0_sel0_signed => x2_2 + to_signed(1,64)
                             , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_0\ ) when \c$~<~Out_case_scrut_2\ else
                             ( Tup2_0_sel0_signed => resPtr_0
                             , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_0\ );

  clash_internal_cOut_0 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_0\
      , xs           => currRes_0
      , ds           => \c$~<~Out_app_arg_2\ );

  \c$~<~Out_app_arg_2\ <= ( Tup2_sel0_signed => x2_2 + to_signed(1,64)
                          , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_0)
                           & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_2\ else
                          \c$~<~Out_case_alt\;

  x2_2 <= resPtr_0;

  with (\c$~<~Out_case_scrut_1\(128 downto 128)) select
    \c$~<~Out_case_alt\ <= ( Tup2_sel0_signed => resPtr_0
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_1)
                            & std_logic_vector(to_signed(1,64))))) ) when "0",
                           ( Tup2_sel0_signed => resPtr_0
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_1)
                            & std_logic_vector(x2_3 + to_signed(1,64))))) ) when others;

  x2_3 <= y_1;

  y_1 <= a1.Tup2_1_sel1_signed_1;

  a1 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_1\(127 downto 0)));

  -- index begin
  indexVec_1 : block
    signal vec_index_1 : integer range 0 to 64-1;
  begin
    vec_index_1 <= to_integer(resPtr_0)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_1\ <= currRes_0(vec_index_1);
  end block;
  -- index end

  currRes_0 <= \c$countConOut_app_arg_0\.Tup2_0_sel1_array_of_Maybe;

  resPtr_0 <= \c$countConOut_app_arg_0\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_2\ <= tagToEnum(\c$~<~Out_app_arg_3\);

  \c$~<~Out_app_arg_3\ <= to_signed(1,64) when x1_0 /= y_2 else to_signed(0,64);

  y_2 <= wild2_1;

  x1_0 <= wild2_0;

  -- index begin
  indexVec_2 : block
    signal vec_index_2 : integer range 0 to 64-1;
  begin
    vec_index_2 <= to_integer(to_signed(62,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_0 <= \c$app_arg\(vec_index_2);
  end block;
  -- index end

  \c$countConOut_app_arg_0\ <= ( Tup2_0_sel0_signed => x2_4 + to_signed(1,64)
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_1\ ) when \c$~<~Out_case_scrut_4\ else
                               ( Tup2_0_sel0_signed => resPtr_1
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_1\ );

  clash_internal_cOut_1 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_1\
      , xs           => currRes_1
      , ds           => \c$~<~Out_app_arg_4\ );

  \c$~<~Out_app_arg_4\ <= ( Tup2_sel0_signed => x2_4 + to_signed(1,64)
                          , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_1)
                           & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_4\ else
                          \c$~<~Out_case_alt_0\;

  x2_4 <= resPtr_1;

  with (\c$~<~Out_case_scrut_3\(128 downto 128)) select
    \c$~<~Out_case_alt_0\ <= ( Tup2_sel0_signed => resPtr_1
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_2)
                              & std_logic_vector(to_signed(1,64))))) ) when "0",
                             ( Tup2_sel0_signed => resPtr_1
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_2)
                              & std_logic_vector(x2_5 + to_signed(1,64))))) ) when others;

  x2_5 <= y_3;

  y_3 <= a1_0.Tup2_1_sel1_signed_1;

  a1_0 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_3\(127 downto 0)));

  -- index begin
  indexVec_3 : block
    signal vec_index_3 : integer range 0 to 64-1;
  begin
    vec_index_3 <= to_integer(resPtr_1)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_3\ <= currRes_1(vec_index_3);
  end block;
  -- index end

  currRes_1 <= \c$countConOut_app_arg_1\.Tup2_0_sel1_array_of_Maybe;

  resPtr_1 <= \c$countConOut_app_arg_1\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_4\ <= tagToEnum(\c$~<~Out_app_arg_5\);

  \c$~<~Out_app_arg_5\ <= to_signed(1,64) when x1_1 /= y_4 else to_signed(0,64);

  y_4 <= wild2_2;

  x1_1 <= wild2_1;

  -- index begin
  indexVec_4 : block
    signal vec_index_4 : integer range 0 to 64-1;
  begin
    vec_index_4 <= to_integer(to_signed(61,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_1 <= \c$app_arg\(vec_index_4);
  end block;
  -- index end

  \c$countConOut_app_arg_1\ <= ( Tup2_0_sel0_signed => x2_6 + to_signed(1,64)
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_2\ ) when \c$~<~Out_case_scrut_6\ else
                               ( Tup2_0_sel0_signed => resPtr_2
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_2\ );

  clash_internal_cOut_2 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_2\
      , xs           => currRes_2
      , ds           => \c$~<~Out_app_arg_6\ );

  \c$~<~Out_app_arg_6\ <= ( Tup2_sel0_signed => x2_6 + to_signed(1,64)
                          , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_2)
                           & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_6\ else
                          \c$~<~Out_case_alt_1\;

  x2_6 <= resPtr_2;

  with (\c$~<~Out_case_scrut_5\(128 downto 128)) select
    \c$~<~Out_case_alt_1\ <= ( Tup2_sel0_signed => resPtr_2
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_3)
                              & std_logic_vector(to_signed(1,64))))) ) when "0",
                             ( Tup2_sel0_signed => resPtr_2
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_3)
                              & std_logic_vector(x2_7 + to_signed(1,64))))) ) when others;

  x2_7 <= y_5;

  y_5 <= a1_1.Tup2_1_sel1_signed_1;

  a1_1 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_5\(127 downto 0)));

  -- index begin
  indexVec_5 : block
    signal vec_index_5 : integer range 0 to 64-1;
  begin
    vec_index_5 <= to_integer(resPtr_2)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_5\ <= currRes_2(vec_index_5);
  end block;
  -- index end

  currRes_2 <= \c$countConOut_app_arg_2\.Tup2_0_sel1_array_of_Maybe;

  resPtr_2 <= \c$countConOut_app_arg_2\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_6\ <= tagToEnum(\c$~<~Out_app_arg_7\);

  \c$~<~Out_app_arg_7\ <= to_signed(1,64) when x1_2 /= y_6 else to_signed(0,64);

  y_6 <= wild2_3;

  x1_2 <= wild2_2;

  -- index begin
  indexVec_6 : block
    signal vec_index_6 : integer range 0 to 64-1;
  begin
    vec_index_6 <= to_integer(to_signed(60,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_2 <= \c$app_arg\(vec_index_6);
  end block;
  -- index end

  \c$countConOut_app_arg_2\ <= ( Tup2_0_sel0_signed => x2_8 + to_signed(1,64)
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_3\ ) when \c$~<~Out_case_scrut_8\ else
                               ( Tup2_0_sel0_signed => resPtr_3
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_3\ );

  clash_internal_cOut_3 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_3\
      , xs           => currRes_3
      , ds           => \c$~<~Out_app_arg_8\ );

  \c$~<~Out_app_arg_8\ <= ( Tup2_sel0_signed => x2_8 + to_signed(1,64)
                          , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_3)
                           & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_8\ else
                          \c$~<~Out_case_alt_2\;

  x2_8 <= resPtr_3;

  with (\c$~<~Out_case_scrut_7\(128 downto 128)) select
    \c$~<~Out_case_alt_2\ <= ( Tup2_sel0_signed => resPtr_3
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_4)
                              & std_logic_vector(to_signed(1,64))))) ) when "0",
                             ( Tup2_sel0_signed => resPtr_3
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_4)
                              & std_logic_vector(x2_9 + to_signed(1,64))))) ) when others;

  x2_9 <= y_7;

  y_7 <= a1_2.Tup2_1_sel1_signed_1;

  a1_2 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_7\(127 downto 0)));

  -- index begin
  indexVec_7 : block
    signal vec_index_7 : integer range 0 to 64-1;
  begin
    vec_index_7 <= to_integer(resPtr_3)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_7\ <= currRes_3(vec_index_7);
  end block;
  -- index end

  currRes_3 <= \c$countConOut_app_arg_3\.Tup2_0_sel1_array_of_Maybe;

  resPtr_3 <= \c$countConOut_app_arg_3\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_8\ <= tagToEnum(\c$~<~Out_app_arg_9\);

  \c$~<~Out_app_arg_9\ <= to_signed(1,64) when x1_3 /= y_8 else to_signed(0,64);

  y_8 <= wild2_4;

  x1_3 <= wild2_3;

  -- index begin
  indexVec_8 : block
    signal vec_index_8 : integer range 0 to 64-1;
  begin
    vec_index_8 <= to_integer(to_signed(59,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_3 <= \c$app_arg\(vec_index_8);
  end block;
  -- index end

  \c$countConOut_app_arg_3\ <= ( Tup2_0_sel0_signed => x2_10 + to_signed(1,64)
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_4\ ) when \c$~<~Out_case_scrut_10\ else
                               ( Tup2_0_sel0_signed => resPtr_4
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_4\ );

  clash_internal_cOut_4 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_4\
      , xs           => currRes_4
      , ds           => \c$~<~Out_app_arg_10\ );

  \c$~<~Out_app_arg_10\ <= ( Tup2_sel0_signed => x2_10 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_4)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_10\ else
                           \c$~<~Out_case_alt_3\;

  x2_10 <= resPtr_4;

  with (\c$~<~Out_case_scrut_9\(128 downto 128)) select
    \c$~<~Out_case_alt_3\ <= ( Tup2_sel0_signed => resPtr_4
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_5)
                              & std_logic_vector(to_signed(1,64))))) ) when "0",
                             ( Tup2_sel0_signed => resPtr_4
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_5)
                              & std_logic_vector(x2_11 + to_signed(1,64))))) ) when others;

  x2_11 <= y_9;

  y_9 <= a1_3.Tup2_1_sel1_signed_1;

  a1_3 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_9\(127 downto 0)));

  -- index begin
  indexVec_9 : block
    signal vec_index_9 : integer range 0 to 64-1;
  begin
    vec_index_9 <= to_integer(resPtr_4)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_9\ <= currRes_4(vec_index_9);
  end block;
  -- index end

  currRes_4 <= \c$countConOut_app_arg_4\.Tup2_0_sel1_array_of_Maybe;

  resPtr_4 <= \c$countConOut_app_arg_4\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_10\ <= tagToEnum(\c$~<~Out_app_arg_11\);

  \c$~<~Out_app_arg_11\ <= to_signed(1,64) when x1_4 /= y_10 else to_signed(0,64);

  y_10 <= wild2_5;

  x1_4 <= wild2_4;

  -- index begin
  indexVec_10 : block
    signal vec_index_10 : integer range 0 to 64-1;
  begin
    vec_index_10 <= to_integer(to_signed(58,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_4 <= \c$app_arg\(vec_index_10);
  end block;
  -- index end

  \c$countConOut_app_arg_4\ <= ( Tup2_0_sel0_signed => x2_12 + to_signed(1,64)
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_5\ ) when \c$~<~Out_case_scrut_12\ else
                               ( Tup2_0_sel0_signed => resPtr_5
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_5\ );

  clash_internal_cOut_5 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_5\
      , xs           => currRes_5
      , ds           => \c$~<~Out_app_arg_12\ );

  \c$~<~Out_app_arg_12\ <= ( Tup2_sel0_signed => x2_12 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_5)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_12\ else
                           \c$~<~Out_case_alt_4\;

  x2_12 <= resPtr_5;

  with (\c$~<~Out_case_scrut_11\(128 downto 128)) select
    \c$~<~Out_case_alt_4\ <= ( Tup2_sel0_signed => resPtr_5
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_6)
                              & std_logic_vector(to_signed(1,64))))) ) when "0",
                             ( Tup2_sel0_signed => resPtr_5
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_6)
                              & std_logic_vector(x2_13 + to_signed(1,64))))) ) when others;

  x2_13 <= y_11;

  y_11 <= a1_4.Tup2_1_sel1_signed_1;

  a1_4 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_11\(127 downto 0)));

  -- index begin
  indexVec_11 : block
    signal vec_index_11 : integer range 0 to 64-1;
  begin
    vec_index_11 <= to_integer(resPtr_5)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_11\ <= currRes_5(vec_index_11);
  end block;
  -- index end

  currRes_5 <= \c$countConOut_app_arg_5\.Tup2_0_sel1_array_of_Maybe;

  resPtr_5 <= \c$countConOut_app_arg_5\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_12\ <= tagToEnum(\c$~<~Out_app_arg_13\);

  \c$~<~Out_app_arg_13\ <= to_signed(1,64) when x1_5 /= y_12 else to_signed(0,64);

  y_12 <= wild2_6;

  x1_5 <= wild2_5;

  -- index begin
  indexVec_12 : block
    signal vec_index_12 : integer range 0 to 64-1;
  begin
    vec_index_12 <= to_integer(to_signed(57,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_5 <= \c$app_arg\(vec_index_12);
  end block;
  -- index end

  \c$countConOut_app_arg_5\ <= ( Tup2_0_sel0_signed => x2_14 + to_signed(1,64)
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_6\ ) when \c$~<~Out_case_scrut_14\ else
                               ( Tup2_0_sel0_signed => resPtr_6
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_6\ );

  clash_internal_cOut_6 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_6\
      , xs           => currRes_6
      , ds           => \c$~<~Out_app_arg_14\ );

  \c$~<~Out_app_arg_14\ <= ( Tup2_sel0_signed => x2_14 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_6)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_14\ else
                           \c$~<~Out_case_alt_5\;

  x2_14 <= resPtr_6;

  with (\c$~<~Out_case_scrut_13\(128 downto 128)) select
    \c$~<~Out_case_alt_5\ <= ( Tup2_sel0_signed => resPtr_6
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_7)
                              & std_logic_vector(to_signed(1,64))))) ) when "0",
                             ( Tup2_sel0_signed => resPtr_6
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_7)
                              & std_logic_vector(x2_15 + to_signed(1,64))))) ) when others;

  x2_15 <= y_13;

  y_13 <= a1_5.Tup2_1_sel1_signed_1;

  a1_5 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_13\(127 downto 0)));

  -- index begin
  indexVec_13 : block
    signal vec_index_13 : integer range 0 to 64-1;
  begin
    vec_index_13 <= to_integer(resPtr_6)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_13\ <= currRes_6(vec_index_13);
  end block;
  -- index end

  currRes_6 <= \c$countConOut_app_arg_6\.Tup2_0_sel1_array_of_Maybe;

  resPtr_6 <= \c$countConOut_app_arg_6\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_14\ <= tagToEnum(\c$~<~Out_app_arg_15\);

  \c$~<~Out_app_arg_15\ <= to_signed(1,64) when x1_6 /= y_14 else to_signed(0,64);

  y_14 <= wild2_7;

  x1_6 <= wild2_6;

  -- index begin
  indexVec_14 : block
    signal vec_index_14 : integer range 0 to 64-1;
  begin
    vec_index_14 <= to_integer(to_signed(56,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_6 <= \c$app_arg\(vec_index_14);
  end block;
  -- index end

  \c$countConOut_app_arg_6\ <= ( Tup2_0_sel0_signed => x2_16 + to_signed(1,64)
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_7\ ) when \c$~<~Out_case_scrut_16\ else
                               ( Tup2_0_sel0_signed => resPtr_7
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_7\ );

  clash_internal_cOut_7 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_7\
      , xs           => currRes_7
      , ds           => \c$~<~Out_app_arg_16\ );

  \c$~<~Out_app_arg_16\ <= ( Tup2_sel0_signed => x2_16 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_7)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_16\ else
                           \c$~<~Out_case_alt_6\;

  x2_16 <= resPtr_7;

  with (\c$~<~Out_case_scrut_15\(128 downto 128)) select
    \c$~<~Out_case_alt_6\ <= ( Tup2_sel0_signed => resPtr_7
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_8)
                              & std_logic_vector(to_signed(1,64))))) ) when "0",
                             ( Tup2_sel0_signed => resPtr_7
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_8)
                              & std_logic_vector(x2_17 + to_signed(1,64))))) ) when others;

  x2_17 <= y_15;

  y_15 <= a1_6.Tup2_1_sel1_signed_1;

  a1_6 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_15\(127 downto 0)));

  -- index begin
  indexVec_15 : block
    signal vec_index_15 : integer range 0 to 64-1;
  begin
    vec_index_15 <= to_integer(resPtr_7)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_15\ <= currRes_7(vec_index_15);
  end block;
  -- index end

  currRes_7 <= \c$countConOut_app_arg_7\.Tup2_0_sel1_array_of_Maybe;

  resPtr_7 <= \c$countConOut_app_arg_7\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_16\ <= tagToEnum(\c$~<~Out_app_arg_17\);

  \c$~<~Out_app_arg_17\ <= to_signed(1,64) when x1_7 /= y_16 else to_signed(0,64);

  y_16 <= wild2_8;

  x1_7 <= wild2_7;

  -- index begin
  indexVec_16 : block
    signal vec_index_16 : integer range 0 to 64-1;
  begin
    vec_index_16 <= to_integer(to_signed(55,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_7 <= \c$app_arg\(vec_index_16);
  end block;
  -- index end

  \c$countConOut_app_arg_7\ <= ( Tup2_0_sel0_signed => x2_18 + to_signed(1,64)
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_8\ ) when \c$~<~Out_case_scrut_18\ else
                               ( Tup2_0_sel0_signed => resPtr_8
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_8\ );

  clash_internal_cOut_8 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_8\
      , xs           => currRes_8
      , ds           => \c$~<~Out_app_arg_18\ );

  \c$~<~Out_app_arg_18\ <= ( Tup2_sel0_signed => x2_18 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_8)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_18\ else
                           \c$~<~Out_case_alt_7\;

  x2_18 <= resPtr_8;

  with (\c$~<~Out_case_scrut_17\(128 downto 128)) select
    \c$~<~Out_case_alt_7\ <= ( Tup2_sel0_signed => resPtr_8
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_9)
                              & std_logic_vector(to_signed(1,64))))) ) when "0",
                             ( Tup2_sel0_signed => resPtr_8
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_9)
                              & std_logic_vector(x2_19 + to_signed(1,64))))) ) when others;

  x2_19 <= y_17;

  y_17 <= a1_7.Tup2_1_sel1_signed_1;

  a1_7 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_17\(127 downto 0)));

  -- index begin
  indexVec_17 : block
    signal vec_index_17 : integer range 0 to 64-1;
  begin
    vec_index_17 <= to_integer(resPtr_8)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_17\ <= currRes_8(vec_index_17);
  end block;
  -- index end

  currRes_8 <= \c$countConOut_app_arg_8\.Tup2_0_sel1_array_of_Maybe;

  resPtr_8 <= \c$countConOut_app_arg_8\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_18\ <= tagToEnum(\c$~<~Out_app_arg_19\);

  \c$~<~Out_app_arg_19\ <= to_signed(1,64) when x1_8 /= y_18 else to_signed(0,64);

  y_18 <= wild2_9;

  x1_8 <= wild2_8;

  -- index begin
  indexVec_18 : block
    signal vec_index_18 : integer range 0 to 64-1;
  begin
    vec_index_18 <= to_integer(to_signed(54,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_8 <= \c$app_arg\(vec_index_18);
  end block;
  -- index end

  \c$countConOut_app_arg_8\ <= ( Tup2_0_sel0_signed => x2_20 + to_signed(1,64)
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_9\ ) when \c$~<~Out_case_scrut_20\ else
                               ( Tup2_0_sel0_signed => resPtr_9
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_9\ );

  clash_internal_cOut_9 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_9\
      , xs           => currRes_9
      , ds           => \c$~<~Out_app_arg_20\ );

  \c$~<~Out_app_arg_20\ <= ( Tup2_sel0_signed => x2_20 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_9)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_20\ else
                           \c$~<~Out_case_alt_8\;

  x2_20 <= resPtr_9;

  with (\c$~<~Out_case_scrut_19\(128 downto 128)) select
    \c$~<~Out_case_alt_8\ <= ( Tup2_sel0_signed => resPtr_9
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_10)
                              & std_logic_vector(to_signed(1,64))))) ) when "0",
                             ( Tup2_sel0_signed => resPtr_9
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_10)
                              & std_logic_vector(x2_21 + to_signed(1,64))))) ) when others;

  x2_21 <= y_19;

  y_19 <= a1_8.Tup2_1_sel1_signed_1;

  a1_8 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_19\(127 downto 0)));

  -- index begin
  indexVec_19 : block
    signal vec_index_19 : integer range 0 to 64-1;
  begin
    vec_index_19 <= to_integer(resPtr_9)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_19\ <= currRes_9(vec_index_19);
  end block;
  -- index end

  currRes_9 <= \c$countConOut_app_arg_9\.Tup2_0_sel1_array_of_Maybe;

  resPtr_9 <= \c$countConOut_app_arg_9\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_20\ <= tagToEnum(\c$~<~Out_app_arg_21\);

  \c$~<~Out_app_arg_21\ <= to_signed(1,64) when x1_9 /= y_20 else to_signed(0,64);

  y_20 <= wild2_10;

  x1_9 <= wild2_9;

  -- index begin
  indexVec_20 : block
    signal vec_index_20 : integer range 0 to 64-1;
  begin
    vec_index_20 <= to_integer(to_signed(53,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_9 <= \c$app_arg\(vec_index_20);
  end block;
  -- index end

  \c$countConOut_app_arg_9\ <= ( Tup2_0_sel0_signed => x2_22 + to_signed(1,64)
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_10\ ) when \c$~<~Out_case_scrut_22\ else
                               ( Tup2_0_sel0_signed => resPtr_10
                               , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_10\ );

  clash_internal_cOut_10 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_10\
      , xs           => currRes_10
      , ds           => \c$~<~Out_app_arg_22\ );

  \c$~<~Out_app_arg_22\ <= ( Tup2_sel0_signed => x2_22 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_10)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_22\ else
                           \c$~<~Out_case_alt_9\;

  x2_22 <= resPtr_10;

  with (\c$~<~Out_case_scrut_21\(128 downto 128)) select
    \c$~<~Out_case_alt_9\ <= ( Tup2_sel0_signed => resPtr_10
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_11)
                              & std_logic_vector(to_signed(1,64))))) ) when "0",
                             ( Tup2_sel0_signed => resPtr_10
                             , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_11)
                              & std_logic_vector(x2_23 + to_signed(1,64))))) ) when others;

  x2_23 <= y_21;

  y_21 <= a1_9.Tup2_1_sel1_signed_1;

  a1_9 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_21\(127 downto 0)));

  -- index begin
  indexVec_21 : block
    signal vec_index_21 : integer range 0 to 64-1;
  begin
    vec_index_21 <= to_integer(resPtr_10)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_21\ <= currRes_10(vec_index_21);
  end block;
  -- index end

  currRes_10 <= \c$countConOut_app_arg_10\.Tup2_0_sel1_array_of_Maybe;

  resPtr_10 <= \c$countConOut_app_arg_10\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_22\ <= tagToEnum(\c$~<~Out_app_arg_23\);

  \c$~<~Out_app_arg_23\ <= to_signed(1,64) when x1_10 /= y_22 else to_signed(0,64);

  y_22 <= wild2_11;

  x1_10 <= wild2_10;

  -- index begin
  indexVec_22 : block
    signal vec_index_22 : integer range 0 to 64-1;
  begin
    vec_index_22 <= to_integer(to_signed(52,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_10 <= \c$app_arg\(vec_index_22);
  end block;
  -- index end

  \c$countConOut_app_arg_10\ <= ( Tup2_0_sel0_signed => x2_24 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_11\ ) when \c$~<~Out_case_scrut_24\ else
                                ( Tup2_0_sel0_signed => resPtr_11
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_11\ );

  clash_internal_cOut_11 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_11\
      , xs           => currRes_11
      , ds           => \c$~<~Out_app_arg_24\ );

  \c$~<~Out_app_arg_24\ <= ( Tup2_sel0_signed => x2_24 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_11)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_24\ else
                           \c$~<~Out_case_alt_10\;

  x2_24 <= resPtr_11;

  with (\c$~<~Out_case_scrut_23\(128 downto 128)) select
    \c$~<~Out_case_alt_10\ <= ( Tup2_sel0_signed => resPtr_11
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_12)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_11
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_12)
                               & std_logic_vector(x2_25 + to_signed(1,64))))) ) when others;

  x2_25 <= y_23;

  y_23 <= a1_10.Tup2_1_sel1_signed_1;

  a1_10 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_23\(127 downto 0)));

  -- index begin
  indexVec_23 : block
    signal vec_index_23 : integer range 0 to 64-1;
  begin
    vec_index_23 <= to_integer(resPtr_11)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_23\ <= currRes_11(vec_index_23);
  end block;
  -- index end

  currRes_11 <= \c$countConOut_app_arg_11\.Tup2_0_sel1_array_of_Maybe;

  resPtr_11 <= \c$countConOut_app_arg_11\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_24\ <= tagToEnum(\c$~<~Out_app_arg_25\);

  \c$~<~Out_app_arg_25\ <= to_signed(1,64) when x1_11 /= y_24 else to_signed(0,64);

  y_24 <= wild2_12;

  x1_11 <= wild2_11;

  -- index begin
  indexVec_24 : block
    signal vec_index_24 : integer range 0 to 64-1;
  begin
    vec_index_24 <= to_integer(to_signed(51,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_11 <= \c$app_arg\(vec_index_24);
  end block;
  -- index end

  \c$countConOut_app_arg_11\ <= ( Tup2_0_sel0_signed => x2_26 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_12\ ) when \c$~<~Out_case_scrut_26\ else
                                ( Tup2_0_sel0_signed => resPtr_12
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_12\ );

  clash_internal_cOut_12 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_12\
      , xs           => currRes_12
      , ds           => \c$~<~Out_app_arg_26\ );

  \c$~<~Out_app_arg_26\ <= ( Tup2_sel0_signed => x2_26 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_12)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_26\ else
                           \c$~<~Out_case_alt_11\;

  x2_26 <= resPtr_12;

  with (\c$~<~Out_case_scrut_25\(128 downto 128)) select
    \c$~<~Out_case_alt_11\ <= ( Tup2_sel0_signed => resPtr_12
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_13)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_12
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_13)
                               & std_logic_vector(x2_27 + to_signed(1,64))))) ) when others;

  x2_27 <= y_25;

  y_25 <= a1_11.Tup2_1_sel1_signed_1;

  a1_11 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_25\(127 downto 0)));

  -- index begin
  indexVec_25 : block
    signal vec_index_25 : integer range 0 to 64-1;
  begin
    vec_index_25 <= to_integer(resPtr_12)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_25\ <= currRes_12(vec_index_25);
  end block;
  -- index end

  currRes_12 <= \c$countConOut_app_arg_12\.Tup2_0_sel1_array_of_Maybe;

  resPtr_12 <= \c$countConOut_app_arg_12\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_26\ <= tagToEnum(\c$~<~Out_app_arg_27\);

  \c$~<~Out_app_arg_27\ <= to_signed(1,64) when x1_12 /= y_26 else to_signed(0,64);

  y_26 <= wild2_13;

  x1_12 <= wild2_12;

  -- index begin
  indexVec_26 : block
    signal vec_index_26 : integer range 0 to 64-1;
  begin
    vec_index_26 <= to_integer(to_signed(50,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_12 <= \c$app_arg\(vec_index_26);
  end block;
  -- index end

  \c$countConOut_app_arg_12\ <= ( Tup2_0_sel0_signed => x2_28 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_13\ ) when \c$~<~Out_case_scrut_28\ else
                                ( Tup2_0_sel0_signed => resPtr_13
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_13\ );

  clash_internal_cOut_13 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_13\
      , xs           => currRes_13
      , ds           => \c$~<~Out_app_arg_28\ );

  \c$~<~Out_app_arg_28\ <= ( Tup2_sel0_signed => x2_28 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_13)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_28\ else
                           \c$~<~Out_case_alt_12\;

  x2_28 <= resPtr_13;

  with (\c$~<~Out_case_scrut_27\(128 downto 128)) select
    \c$~<~Out_case_alt_12\ <= ( Tup2_sel0_signed => resPtr_13
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_14)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_13
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_14)
                               & std_logic_vector(x2_29 + to_signed(1,64))))) ) when others;

  x2_29 <= y_27;

  y_27 <= a1_12.Tup2_1_sel1_signed_1;

  a1_12 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_27\(127 downto 0)));

  -- index begin
  indexVec_27 : block
    signal vec_index_27 : integer range 0 to 64-1;
  begin
    vec_index_27 <= to_integer(resPtr_13)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_27\ <= currRes_13(vec_index_27);
  end block;
  -- index end

  currRes_13 <= \c$countConOut_app_arg_13\.Tup2_0_sel1_array_of_Maybe;

  resPtr_13 <= \c$countConOut_app_arg_13\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_28\ <= tagToEnum(\c$~<~Out_app_arg_29\);

  \c$~<~Out_app_arg_29\ <= to_signed(1,64) when x1_13 /= y_28 else to_signed(0,64);

  y_28 <= wild2_14;

  x1_13 <= wild2_13;

  -- index begin
  indexVec_28 : block
    signal vec_index_28 : integer range 0 to 64-1;
  begin
    vec_index_28 <= to_integer(to_signed(49,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_13 <= \c$app_arg\(vec_index_28);
  end block;
  -- index end

  \c$countConOut_app_arg_13\ <= ( Tup2_0_sel0_signed => x2_30 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_14\ ) when \c$~<~Out_case_scrut_30\ else
                                ( Tup2_0_sel0_signed => resPtr_14
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_14\ );

  clash_internal_cOut_14 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_14\
      , xs           => currRes_14
      , ds           => \c$~<~Out_app_arg_30\ );

  \c$~<~Out_app_arg_30\ <= ( Tup2_sel0_signed => x2_30 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_14)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_30\ else
                           \c$~<~Out_case_alt_13\;

  x2_30 <= resPtr_14;

  with (\c$~<~Out_case_scrut_29\(128 downto 128)) select
    \c$~<~Out_case_alt_13\ <= ( Tup2_sel0_signed => resPtr_14
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_15)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_14
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_15)
                               & std_logic_vector(x2_31 + to_signed(1,64))))) ) when others;

  x2_31 <= y_29;

  y_29 <= a1_13.Tup2_1_sel1_signed_1;

  a1_13 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_29\(127 downto 0)));

  -- index begin
  indexVec_29 : block
    signal vec_index_29 : integer range 0 to 64-1;
  begin
    vec_index_29 <= to_integer(resPtr_14)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_29\ <= currRes_14(vec_index_29);
  end block;
  -- index end

  currRes_14 <= \c$countConOut_app_arg_14\.Tup2_0_sel1_array_of_Maybe;

  resPtr_14 <= \c$countConOut_app_arg_14\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_30\ <= tagToEnum(\c$~<~Out_app_arg_31\);

  \c$~<~Out_app_arg_31\ <= to_signed(1,64) when x1_14 /= y_30 else to_signed(0,64);

  y_30 <= wild2_15;

  x1_14 <= wild2_14;

  -- index begin
  indexVec_30 : block
    signal vec_index_30 : integer range 0 to 64-1;
  begin
    vec_index_30 <= to_integer(to_signed(48,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_14 <= \c$app_arg\(vec_index_30);
  end block;
  -- index end

  \c$countConOut_app_arg_14\ <= ( Tup2_0_sel0_signed => x2_32 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_15\ ) when \c$~<~Out_case_scrut_32\ else
                                ( Tup2_0_sel0_signed => resPtr_15
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_15\ );

  clash_internal_cOut_15 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_15\
      , xs           => currRes_15
      , ds           => \c$~<~Out_app_arg_32\ );

  \c$~<~Out_app_arg_32\ <= ( Tup2_sel0_signed => x2_32 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_15)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_32\ else
                           \c$~<~Out_case_alt_14\;

  x2_32 <= resPtr_15;

  with (\c$~<~Out_case_scrut_31\(128 downto 128)) select
    \c$~<~Out_case_alt_14\ <= ( Tup2_sel0_signed => resPtr_15
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_16)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_15
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_16)
                               & std_logic_vector(x2_33 + to_signed(1,64))))) ) when others;

  x2_33 <= y_31;

  y_31 <= a1_14.Tup2_1_sel1_signed_1;

  a1_14 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_31\(127 downto 0)));

  -- index begin
  indexVec_31 : block
    signal vec_index_31 : integer range 0 to 64-1;
  begin
    vec_index_31 <= to_integer(resPtr_15)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_31\ <= currRes_15(vec_index_31);
  end block;
  -- index end

  currRes_15 <= \c$countConOut_app_arg_15\.Tup2_0_sel1_array_of_Maybe;

  resPtr_15 <= \c$countConOut_app_arg_15\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_32\ <= tagToEnum(\c$~<~Out_app_arg_33\);

  \c$~<~Out_app_arg_33\ <= to_signed(1,64) when x1_15 /= y_32 else to_signed(0,64);

  y_32 <= wild2_16;

  x1_15 <= wild2_15;

  -- index begin
  indexVec_32 : block
    signal vec_index_32 : integer range 0 to 64-1;
  begin
    vec_index_32 <= to_integer(to_signed(47,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_15 <= \c$app_arg\(vec_index_32);
  end block;
  -- index end

  \c$countConOut_app_arg_15\ <= ( Tup2_0_sel0_signed => x2_34 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_16\ ) when \c$~<~Out_case_scrut_34\ else
                                ( Tup2_0_sel0_signed => resPtr_16
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_16\ );

  clash_internal_cOut_16 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_16\
      , xs           => currRes_16
      , ds           => \c$~<~Out_app_arg_34\ );

  \c$~<~Out_app_arg_34\ <= ( Tup2_sel0_signed => x2_34 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_16)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_34\ else
                           \c$~<~Out_case_alt_15\;

  x2_34 <= resPtr_16;

  with (\c$~<~Out_case_scrut_33\(128 downto 128)) select
    \c$~<~Out_case_alt_15\ <= ( Tup2_sel0_signed => resPtr_16
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_17)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_16
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_17)
                               & std_logic_vector(x2_35 + to_signed(1,64))))) ) when others;

  x2_35 <= y_33;

  y_33 <= a1_15.Tup2_1_sel1_signed_1;

  a1_15 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_33\(127 downto 0)));

  -- index begin
  indexVec_33 : block
    signal vec_index_33 : integer range 0 to 64-1;
  begin
    vec_index_33 <= to_integer(resPtr_16)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_33\ <= currRes_16(vec_index_33);
  end block;
  -- index end

  currRes_16 <= \c$countConOut_app_arg_16\.Tup2_0_sel1_array_of_Maybe;

  resPtr_16 <= \c$countConOut_app_arg_16\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_34\ <= tagToEnum(\c$~<~Out_app_arg_35\);

  \c$~<~Out_app_arg_35\ <= to_signed(1,64) when x1_16 /= y_34 else to_signed(0,64);

  y_34 <= wild2_17;

  x1_16 <= wild2_16;

  -- index begin
  indexVec_34 : block
    signal vec_index_34 : integer range 0 to 64-1;
  begin
    vec_index_34 <= to_integer(to_signed(46,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_16 <= \c$app_arg\(vec_index_34);
  end block;
  -- index end

  \c$countConOut_app_arg_16\ <= ( Tup2_0_sel0_signed => x2_36 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_17\ ) when \c$~<~Out_case_scrut_36\ else
                                ( Tup2_0_sel0_signed => resPtr_17
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_17\ );

  clash_internal_cOut_17 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_17\
      , xs           => currRes_17
      , ds           => \c$~<~Out_app_arg_36\ );

  \c$~<~Out_app_arg_36\ <= ( Tup2_sel0_signed => x2_36 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_17)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_36\ else
                           \c$~<~Out_case_alt_16\;

  x2_36 <= resPtr_17;

  with (\c$~<~Out_case_scrut_35\(128 downto 128)) select
    \c$~<~Out_case_alt_16\ <= ( Tup2_sel0_signed => resPtr_17
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_18)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_17
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_18)
                               & std_logic_vector(x2_37 + to_signed(1,64))))) ) when others;

  x2_37 <= y_35;

  y_35 <= a1_16.Tup2_1_sel1_signed_1;

  a1_16 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_35\(127 downto 0)));

  -- index begin
  indexVec_35 : block
    signal vec_index_35 : integer range 0 to 64-1;
  begin
    vec_index_35 <= to_integer(resPtr_17)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_35\ <= currRes_17(vec_index_35);
  end block;
  -- index end

  currRes_17 <= \c$countConOut_app_arg_17\.Tup2_0_sel1_array_of_Maybe;

  resPtr_17 <= \c$countConOut_app_arg_17\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_36\ <= tagToEnum(\c$~<~Out_app_arg_37\);

  \c$~<~Out_app_arg_37\ <= to_signed(1,64) when x1_17 /= y_36 else to_signed(0,64);

  y_36 <= wild2_18;

  x1_17 <= wild2_17;

  -- index begin
  indexVec_36 : block
    signal vec_index_36 : integer range 0 to 64-1;
  begin
    vec_index_36 <= to_integer(to_signed(45,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_17 <= \c$app_arg\(vec_index_36);
  end block;
  -- index end

  \c$countConOut_app_arg_17\ <= ( Tup2_0_sel0_signed => x2_38 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_18\ ) when \c$~<~Out_case_scrut_38\ else
                                ( Tup2_0_sel0_signed => resPtr_18
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_18\ );

  clash_internal_cOut_18 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_18\
      , xs           => currRes_18
      , ds           => \c$~<~Out_app_arg_38\ );

  \c$~<~Out_app_arg_38\ <= ( Tup2_sel0_signed => x2_38 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_18)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_38\ else
                           \c$~<~Out_case_alt_17\;

  x2_38 <= resPtr_18;

  with (\c$~<~Out_case_scrut_37\(128 downto 128)) select
    \c$~<~Out_case_alt_17\ <= ( Tup2_sel0_signed => resPtr_18
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_19)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_18
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_19)
                               & std_logic_vector(x2_39 + to_signed(1,64))))) ) when others;

  x2_39 <= y_37;

  y_37 <= a1_17.Tup2_1_sel1_signed_1;

  a1_17 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_37\(127 downto 0)));

  -- index begin
  indexVec_37 : block
    signal vec_index_37 : integer range 0 to 64-1;
  begin
    vec_index_37 <= to_integer(resPtr_18)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_37\ <= currRes_18(vec_index_37);
  end block;
  -- index end

  currRes_18 <= \c$countConOut_app_arg_18\.Tup2_0_sel1_array_of_Maybe;

  resPtr_18 <= \c$countConOut_app_arg_18\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_38\ <= tagToEnum(\c$~<~Out_app_arg_39\);

  \c$~<~Out_app_arg_39\ <= to_signed(1,64) when x1_18 /= y_38 else to_signed(0,64);

  y_38 <= wild2_19;

  x1_18 <= wild2_18;

  -- index begin
  indexVec_38 : block
    signal vec_index_38 : integer range 0 to 64-1;
  begin
    vec_index_38 <= to_integer(to_signed(44,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_18 <= \c$app_arg\(vec_index_38);
  end block;
  -- index end

  \c$countConOut_app_arg_18\ <= ( Tup2_0_sel0_signed => x2_40 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_19\ ) when \c$~<~Out_case_scrut_40\ else
                                ( Tup2_0_sel0_signed => resPtr_19
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_19\ );

  clash_internal_cOut_19 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_19\
      , xs           => currRes_19
      , ds           => \c$~<~Out_app_arg_40\ );

  \c$~<~Out_app_arg_40\ <= ( Tup2_sel0_signed => x2_40 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_19)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_40\ else
                           \c$~<~Out_case_alt_18\;

  x2_40 <= resPtr_19;

  with (\c$~<~Out_case_scrut_39\(128 downto 128)) select
    \c$~<~Out_case_alt_18\ <= ( Tup2_sel0_signed => resPtr_19
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_20)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_19
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_20)
                               & std_logic_vector(x2_41 + to_signed(1,64))))) ) when others;

  x2_41 <= y_39;

  y_39 <= a1_18.Tup2_1_sel1_signed_1;

  a1_18 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_39\(127 downto 0)));

  -- index begin
  indexVec_39 : block
    signal vec_index_39 : integer range 0 to 64-1;
  begin
    vec_index_39 <= to_integer(resPtr_19)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_39\ <= currRes_19(vec_index_39);
  end block;
  -- index end

  currRes_19 <= \c$countConOut_app_arg_19\.Tup2_0_sel1_array_of_Maybe;

  resPtr_19 <= \c$countConOut_app_arg_19\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_40\ <= tagToEnum(\c$~<~Out_app_arg_41\);

  \c$~<~Out_app_arg_41\ <= to_signed(1,64) when x1_19 /= y_40 else to_signed(0,64);

  y_40 <= wild2_20;

  x1_19 <= wild2_19;

  -- index begin
  indexVec_40 : block
    signal vec_index_40 : integer range 0 to 64-1;
  begin
    vec_index_40 <= to_integer(to_signed(43,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_19 <= \c$app_arg\(vec_index_40);
  end block;
  -- index end

  \c$countConOut_app_arg_19\ <= ( Tup2_0_sel0_signed => x2_42 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_20\ ) when \c$~<~Out_case_scrut_42\ else
                                ( Tup2_0_sel0_signed => resPtr_20
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_20\ );

  clash_internal_cOut_20 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_20\
      , xs           => currRes_20
      , ds           => \c$~<~Out_app_arg_42\ );

  \c$~<~Out_app_arg_42\ <= ( Tup2_sel0_signed => x2_42 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_20)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_42\ else
                           \c$~<~Out_case_alt_19\;

  x2_42 <= resPtr_20;

  with (\c$~<~Out_case_scrut_41\(128 downto 128)) select
    \c$~<~Out_case_alt_19\ <= ( Tup2_sel0_signed => resPtr_20
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_21)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_20
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_21)
                               & std_logic_vector(x2_43 + to_signed(1,64))))) ) when others;

  x2_43 <= y_41;

  y_41 <= a1_19.Tup2_1_sel1_signed_1;

  a1_19 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_41\(127 downto 0)));

  -- index begin
  indexVec_41 : block
    signal vec_index_41 : integer range 0 to 64-1;
  begin
    vec_index_41 <= to_integer(resPtr_20)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_41\ <= currRes_20(vec_index_41);
  end block;
  -- index end

  currRes_20 <= \c$countConOut_app_arg_20\.Tup2_0_sel1_array_of_Maybe;

  resPtr_20 <= \c$countConOut_app_arg_20\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_42\ <= tagToEnum(\c$~<~Out_app_arg_43\);

  \c$~<~Out_app_arg_43\ <= to_signed(1,64) when x1_20 /= y_42 else to_signed(0,64);

  y_42 <= wild2_21;

  x1_20 <= wild2_20;

  -- index begin
  indexVec_42 : block
    signal vec_index_42 : integer range 0 to 64-1;
  begin
    vec_index_42 <= to_integer(to_signed(42,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_20 <= \c$app_arg\(vec_index_42);
  end block;
  -- index end

  \c$countConOut_app_arg_20\ <= ( Tup2_0_sel0_signed => x2_44 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_21\ ) when \c$~<~Out_case_scrut_44\ else
                                ( Tup2_0_sel0_signed => resPtr_21
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_21\ );

  clash_internal_cOut_21 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_21\
      , xs           => currRes_21
      , ds           => \c$~<~Out_app_arg_44\ );

  \c$~<~Out_app_arg_44\ <= ( Tup2_sel0_signed => x2_44 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_21)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_44\ else
                           \c$~<~Out_case_alt_20\;

  x2_44 <= resPtr_21;

  with (\c$~<~Out_case_scrut_43\(128 downto 128)) select
    \c$~<~Out_case_alt_20\ <= ( Tup2_sel0_signed => resPtr_21
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_22)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_21
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_22)
                               & std_logic_vector(x2_45 + to_signed(1,64))))) ) when others;

  x2_45 <= y_43;

  y_43 <= a1_20.Tup2_1_sel1_signed_1;

  a1_20 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_43\(127 downto 0)));

  -- index begin
  indexVec_43 : block
    signal vec_index_43 : integer range 0 to 64-1;
  begin
    vec_index_43 <= to_integer(resPtr_21)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_43\ <= currRes_21(vec_index_43);
  end block;
  -- index end

  currRes_21 <= \c$countConOut_app_arg_21\.Tup2_0_sel1_array_of_Maybe;

  resPtr_21 <= \c$countConOut_app_arg_21\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_44\ <= tagToEnum(\c$~<~Out_app_arg_45\);

  \c$~<~Out_app_arg_45\ <= to_signed(1,64) when x1_21 /= y_44 else to_signed(0,64);

  y_44 <= wild2_22;

  x1_21 <= wild2_21;

  -- index begin
  indexVec_44 : block
    signal vec_index_44 : integer range 0 to 64-1;
  begin
    vec_index_44 <= to_integer(to_signed(41,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_21 <= \c$app_arg\(vec_index_44);
  end block;
  -- index end

  \c$countConOut_app_arg_21\ <= ( Tup2_0_sel0_signed => x2_46 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_22\ ) when \c$~<~Out_case_scrut_46\ else
                                ( Tup2_0_sel0_signed => resPtr_22
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_22\ );

  clash_internal_cOut_22 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_22\
      , xs           => currRes_22
      , ds           => \c$~<~Out_app_arg_46\ );

  \c$~<~Out_app_arg_46\ <= ( Tup2_sel0_signed => x2_46 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_22)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_46\ else
                           \c$~<~Out_case_alt_21\;

  x2_46 <= resPtr_22;

  with (\c$~<~Out_case_scrut_45\(128 downto 128)) select
    \c$~<~Out_case_alt_21\ <= ( Tup2_sel0_signed => resPtr_22
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_23)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_22
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_23)
                               & std_logic_vector(x2_47 + to_signed(1,64))))) ) when others;

  x2_47 <= y_45;

  y_45 <= a1_21.Tup2_1_sel1_signed_1;

  a1_21 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_45\(127 downto 0)));

  -- index begin
  indexVec_45 : block
    signal vec_index_45 : integer range 0 to 64-1;
  begin
    vec_index_45 <= to_integer(resPtr_22)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_45\ <= currRes_22(vec_index_45);
  end block;
  -- index end

  currRes_22 <= \c$countConOut_app_arg_22\.Tup2_0_sel1_array_of_Maybe;

  resPtr_22 <= \c$countConOut_app_arg_22\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_46\ <= tagToEnum(\c$~<~Out_app_arg_47\);

  \c$~<~Out_app_arg_47\ <= to_signed(1,64) when x1_22 /= y_46 else to_signed(0,64);

  y_46 <= wild2_23;

  x1_22 <= wild2_22;

  -- index begin
  indexVec_46 : block
    signal vec_index_46 : integer range 0 to 64-1;
  begin
    vec_index_46 <= to_integer(to_signed(40,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_22 <= \c$app_arg\(vec_index_46);
  end block;
  -- index end

  \c$countConOut_app_arg_22\ <= ( Tup2_0_sel0_signed => x2_48 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_23\ ) when \c$~<~Out_case_scrut_48\ else
                                ( Tup2_0_sel0_signed => resPtr_23
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_23\ );

  clash_internal_cOut_23 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_23\
      , xs           => currRes_23
      , ds           => \c$~<~Out_app_arg_48\ );

  \c$~<~Out_app_arg_48\ <= ( Tup2_sel0_signed => x2_48 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_23)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_48\ else
                           \c$~<~Out_case_alt_22\;

  x2_48 <= resPtr_23;

  with (\c$~<~Out_case_scrut_47\(128 downto 128)) select
    \c$~<~Out_case_alt_22\ <= ( Tup2_sel0_signed => resPtr_23
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_24)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_23
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_24)
                               & std_logic_vector(x2_49 + to_signed(1,64))))) ) when others;

  x2_49 <= y_47;

  y_47 <= a1_22.Tup2_1_sel1_signed_1;

  a1_22 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_47\(127 downto 0)));

  -- index begin
  indexVec_47 : block
    signal vec_index_47 : integer range 0 to 64-1;
  begin
    vec_index_47 <= to_integer(resPtr_23)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_47\ <= currRes_23(vec_index_47);
  end block;
  -- index end

  currRes_23 <= \c$countConOut_app_arg_23\.Tup2_0_sel1_array_of_Maybe;

  resPtr_23 <= \c$countConOut_app_arg_23\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_48\ <= tagToEnum(\c$~<~Out_app_arg_49\);

  \c$~<~Out_app_arg_49\ <= to_signed(1,64) when x1_23 /= y_48 else to_signed(0,64);

  y_48 <= wild2_24;

  x1_23 <= wild2_23;

  -- index begin
  indexVec_48 : block
    signal vec_index_48 : integer range 0 to 64-1;
  begin
    vec_index_48 <= to_integer(to_signed(39,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_23 <= \c$app_arg\(vec_index_48);
  end block;
  -- index end

  \c$countConOut_app_arg_23\ <= ( Tup2_0_sel0_signed => x2_50 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_24\ ) when \c$~<~Out_case_scrut_50\ else
                                ( Tup2_0_sel0_signed => resPtr_24
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_24\ );

  clash_internal_cOut_24 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_24\
      , xs           => currRes_24
      , ds           => \c$~<~Out_app_arg_50\ );

  \c$~<~Out_app_arg_50\ <= ( Tup2_sel0_signed => x2_50 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_24)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_50\ else
                           \c$~<~Out_case_alt_23\;

  x2_50 <= resPtr_24;

  with (\c$~<~Out_case_scrut_49\(128 downto 128)) select
    \c$~<~Out_case_alt_23\ <= ( Tup2_sel0_signed => resPtr_24
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_25)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_24
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_25)
                               & std_logic_vector(x2_51 + to_signed(1,64))))) ) when others;

  x2_51 <= y_49;

  y_49 <= a1_23.Tup2_1_sel1_signed_1;

  a1_23 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_49\(127 downto 0)));

  -- index begin
  indexVec_49 : block
    signal vec_index_49 : integer range 0 to 64-1;
  begin
    vec_index_49 <= to_integer(resPtr_24)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_49\ <= currRes_24(vec_index_49);
  end block;
  -- index end

  currRes_24 <= \c$countConOut_app_arg_24\.Tup2_0_sel1_array_of_Maybe;

  resPtr_24 <= \c$countConOut_app_arg_24\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_50\ <= tagToEnum(\c$~<~Out_app_arg_51\);

  \c$~<~Out_app_arg_51\ <= to_signed(1,64) when x1_24 /= y_50 else to_signed(0,64);

  y_50 <= wild2_25;

  x1_24 <= wild2_24;

  -- index begin
  indexVec_50 : block
    signal vec_index_50 : integer range 0 to 64-1;
  begin
    vec_index_50 <= to_integer(to_signed(38,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_24 <= \c$app_arg\(vec_index_50);
  end block;
  -- index end

  \c$countConOut_app_arg_24\ <= ( Tup2_0_sel0_signed => x2_52 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_25\ ) when \c$~<~Out_case_scrut_52\ else
                                ( Tup2_0_sel0_signed => resPtr_25
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_25\ );

  clash_internal_cOut_25 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_25\
      , xs           => currRes_25
      , ds           => \c$~<~Out_app_arg_52\ );

  \c$~<~Out_app_arg_52\ <= ( Tup2_sel0_signed => x2_52 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_25)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_52\ else
                           \c$~<~Out_case_alt_24\;

  x2_52 <= resPtr_25;

  with (\c$~<~Out_case_scrut_51\(128 downto 128)) select
    \c$~<~Out_case_alt_24\ <= ( Tup2_sel0_signed => resPtr_25
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_26)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_25
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_26)
                               & std_logic_vector(x2_53 + to_signed(1,64))))) ) when others;

  x2_53 <= y_51;

  y_51 <= a1_24.Tup2_1_sel1_signed_1;

  a1_24 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_51\(127 downto 0)));

  -- index begin
  indexVec_51 : block
    signal vec_index_51 : integer range 0 to 64-1;
  begin
    vec_index_51 <= to_integer(resPtr_25)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_51\ <= currRes_25(vec_index_51);
  end block;
  -- index end

  currRes_25 <= \c$countConOut_app_arg_25\.Tup2_0_sel1_array_of_Maybe;

  resPtr_25 <= \c$countConOut_app_arg_25\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_52\ <= tagToEnum(\c$~<~Out_app_arg_53\);

  \c$~<~Out_app_arg_53\ <= to_signed(1,64) when x1_25 /= y_52 else to_signed(0,64);

  y_52 <= wild2_26;

  x1_25 <= wild2_25;

  -- index begin
  indexVec_52 : block
    signal vec_index_52 : integer range 0 to 64-1;
  begin
    vec_index_52 <= to_integer(to_signed(37,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_25 <= \c$app_arg\(vec_index_52);
  end block;
  -- index end

  \c$countConOut_app_arg_25\ <= ( Tup2_0_sel0_signed => x2_54 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_26\ ) when \c$~<~Out_case_scrut_54\ else
                                ( Tup2_0_sel0_signed => resPtr_26
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_26\ );

  clash_internal_cOut_26 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_26\
      , xs           => currRes_26
      , ds           => \c$~<~Out_app_arg_54\ );

  \c$~<~Out_app_arg_54\ <= ( Tup2_sel0_signed => x2_54 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_26)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_54\ else
                           \c$~<~Out_case_alt_25\;

  x2_54 <= resPtr_26;

  with (\c$~<~Out_case_scrut_53\(128 downto 128)) select
    \c$~<~Out_case_alt_25\ <= ( Tup2_sel0_signed => resPtr_26
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_27)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_26
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_27)
                               & std_logic_vector(x2_55 + to_signed(1,64))))) ) when others;

  x2_55 <= y_53;

  y_53 <= a1_25.Tup2_1_sel1_signed_1;

  a1_25 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_53\(127 downto 0)));

  -- index begin
  indexVec_53 : block
    signal vec_index_53 : integer range 0 to 64-1;
  begin
    vec_index_53 <= to_integer(resPtr_26)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_53\ <= currRes_26(vec_index_53);
  end block;
  -- index end

  currRes_26 <= \c$countConOut_app_arg_26\.Tup2_0_sel1_array_of_Maybe;

  resPtr_26 <= \c$countConOut_app_arg_26\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_54\ <= tagToEnum(\c$~<~Out_app_arg_55\);

  \c$~<~Out_app_arg_55\ <= to_signed(1,64) when x1_26 /= y_54 else to_signed(0,64);

  y_54 <= wild2_27;

  x1_26 <= wild2_26;

  -- index begin
  indexVec_54 : block
    signal vec_index_54 : integer range 0 to 64-1;
  begin
    vec_index_54 <= to_integer(to_signed(36,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_26 <= \c$app_arg\(vec_index_54);
  end block;
  -- index end

  \c$countConOut_app_arg_26\ <= ( Tup2_0_sel0_signed => x2_56 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_27\ ) when \c$~<~Out_case_scrut_56\ else
                                ( Tup2_0_sel0_signed => resPtr_27
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_27\ );

  clash_internal_cOut_27 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_27\
      , xs           => currRes_27
      , ds           => \c$~<~Out_app_arg_56\ );

  \c$~<~Out_app_arg_56\ <= ( Tup2_sel0_signed => x2_56 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_27)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_56\ else
                           \c$~<~Out_case_alt_26\;

  x2_56 <= resPtr_27;

  with (\c$~<~Out_case_scrut_55\(128 downto 128)) select
    \c$~<~Out_case_alt_26\ <= ( Tup2_sel0_signed => resPtr_27
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_28)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_27
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_28)
                               & std_logic_vector(x2_57 + to_signed(1,64))))) ) when others;

  x2_57 <= y_55;

  y_55 <= a1_26.Tup2_1_sel1_signed_1;

  a1_26 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_55\(127 downto 0)));

  -- index begin
  indexVec_55 : block
    signal vec_index_55 : integer range 0 to 64-1;
  begin
    vec_index_55 <= to_integer(resPtr_27)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_55\ <= currRes_27(vec_index_55);
  end block;
  -- index end

  currRes_27 <= \c$countConOut_app_arg_27\.Tup2_0_sel1_array_of_Maybe;

  resPtr_27 <= \c$countConOut_app_arg_27\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_56\ <= tagToEnum(\c$~<~Out_app_arg_57\);

  \c$~<~Out_app_arg_57\ <= to_signed(1,64) when x1_27 /= y_56 else to_signed(0,64);

  y_56 <= wild2_28;

  x1_27 <= wild2_27;

  -- index begin
  indexVec_56 : block
    signal vec_index_56 : integer range 0 to 64-1;
  begin
    vec_index_56 <= to_integer(to_signed(35,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_27 <= \c$app_arg\(vec_index_56);
  end block;
  -- index end

  \c$countConOut_app_arg_27\ <= ( Tup2_0_sel0_signed => x2_58 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_28\ ) when \c$~<~Out_case_scrut_58\ else
                                ( Tup2_0_sel0_signed => resPtr_28
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_28\ );

  clash_internal_cOut_28 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_28\
      , xs           => currRes_28
      , ds           => \c$~<~Out_app_arg_58\ );

  \c$~<~Out_app_arg_58\ <= ( Tup2_sel0_signed => x2_58 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_28)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_58\ else
                           \c$~<~Out_case_alt_27\;

  x2_58 <= resPtr_28;

  with (\c$~<~Out_case_scrut_57\(128 downto 128)) select
    \c$~<~Out_case_alt_27\ <= ( Tup2_sel0_signed => resPtr_28
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_29)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_28
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_29)
                               & std_logic_vector(x2_59 + to_signed(1,64))))) ) when others;

  x2_59 <= y_57;

  y_57 <= a1_27.Tup2_1_sel1_signed_1;

  a1_27 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_57\(127 downto 0)));

  -- index begin
  indexVec_57 : block
    signal vec_index_57 : integer range 0 to 64-1;
  begin
    vec_index_57 <= to_integer(resPtr_28)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_57\ <= currRes_28(vec_index_57);
  end block;
  -- index end

  currRes_28 <= \c$countConOut_app_arg_28\.Tup2_0_sel1_array_of_Maybe;

  resPtr_28 <= \c$countConOut_app_arg_28\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_58\ <= tagToEnum(\c$~<~Out_app_arg_59\);

  \c$~<~Out_app_arg_59\ <= to_signed(1,64) when x1_28 /= y_58 else to_signed(0,64);

  y_58 <= wild2_29;

  x1_28 <= wild2_28;

  -- index begin
  indexVec_58 : block
    signal vec_index_58 : integer range 0 to 64-1;
  begin
    vec_index_58 <= to_integer(to_signed(34,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_28 <= \c$app_arg\(vec_index_58);
  end block;
  -- index end

  \c$countConOut_app_arg_28\ <= ( Tup2_0_sel0_signed => x2_60 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_29\ ) when \c$~<~Out_case_scrut_60\ else
                                ( Tup2_0_sel0_signed => resPtr_29
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_29\ );

  clash_internal_cOut_29 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_29\
      , xs           => currRes_29
      , ds           => \c$~<~Out_app_arg_60\ );

  \c$~<~Out_app_arg_60\ <= ( Tup2_sel0_signed => x2_60 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_29)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_60\ else
                           \c$~<~Out_case_alt_28\;

  x2_60 <= resPtr_29;

  with (\c$~<~Out_case_scrut_59\(128 downto 128)) select
    \c$~<~Out_case_alt_28\ <= ( Tup2_sel0_signed => resPtr_29
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_30)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_29
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_30)
                               & std_logic_vector(x2_61 + to_signed(1,64))))) ) when others;

  x2_61 <= y_59;

  y_59 <= a1_28.Tup2_1_sel1_signed_1;

  a1_28 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_59\(127 downto 0)));

  -- index begin
  indexVec_59 : block
    signal vec_index_59 : integer range 0 to 64-1;
  begin
    vec_index_59 <= to_integer(resPtr_29)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_59\ <= currRes_29(vec_index_59);
  end block;
  -- index end

  currRes_29 <= \c$countConOut_app_arg_29\.Tup2_0_sel1_array_of_Maybe;

  resPtr_29 <= \c$countConOut_app_arg_29\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_60\ <= tagToEnum(\c$~<~Out_app_arg_61\);

  \c$~<~Out_app_arg_61\ <= to_signed(1,64) when x1_29 /= y_60 else to_signed(0,64);

  y_60 <= wild2_30;

  x1_29 <= wild2_29;

  -- index begin
  indexVec_60 : block
    signal vec_index_60 : integer range 0 to 64-1;
  begin
    vec_index_60 <= to_integer(to_signed(33,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_29 <= \c$app_arg\(vec_index_60);
  end block;
  -- index end

  \c$countConOut_app_arg_29\ <= ( Tup2_0_sel0_signed => x2_62 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_30\ ) when \c$~<~Out_case_scrut_62\ else
                                ( Tup2_0_sel0_signed => resPtr_30
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_30\ );

  clash_internal_cOut_30 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_30\
      , xs           => currRes_30
      , ds           => \c$~<~Out_app_arg_62\ );

  \c$~<~Out_app_arg_62\ <= ( Tup2_sel0_signed => x2_62 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_30)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_62\ else
                           \c$~<~Out_case_alt_29\;

  x2_62 <= resPtr_30;

  with (\c$~<~Out_case_scrut_61\(128 downto 128)) select
    \c$~<~Out_case_alt_29\ <= ( Tup2_sel0_signed => resPtr_30
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_31)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_30
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_31)
                               & std_logic_vector(x2_63 + to_signed(1,64))))) ) when others;

  x2_63 <= y_61;

  y_61 <= a1_29.Tup2_1_sel1_signed_1;

  a1_29 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_61\(127 downto 0)));

  -- index begin
  indexVec_61 : block
    signal vec_index_61 : integer range 0 to 64-1;
  begin
    vec_index_61 <= to_integer(resPtr_30)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_61\ <= currRes_30(vec_index_61);
  end block;
  -- index end

  currRes_30 <= \c$countConOut_app_arg_30\.Tup2_0_sel1_array_of_Maybe;

  resPtr_30 <= \c$countConOut_app_arg_30\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_62\ <= tagToEnum(\c$~<~Out_app_arg_63\);

  \c$~<~Out_app_arg_63\ <= to_signed(1,64) when x1_30 /= y_62 else to_signed(0,64);

  y_62 <= wild2_31;

  x1_30 <= wild2_30;

  -- index begin
  indexVec_62 : block
    signal vec_index_62 : integer range 0 to 64-1;
  begin
    vec_index_62 <= to_integer(to_signed(32,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_30 <= \c$app_arg\(vec_index_62);
  end block;
  -- index end

  \c$countConOut_app_arg_30\ <= ( Tup2_0_sel0_signed => x2_64 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_31\ ) when \c$~<~Out_case_scrut_64\ else
                                ( Tup2_0_sel0_signed => resPtr_31
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_31\ );

  clash_internal_cOut_31 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_31\
      , xs           => currRes_31
      , ds           => \c$~<~Out_app_arg_64\ );

  \c$~<~Out_app_arg_64\ <= ( Tup2_sel0_signed => x2_64 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_31)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_64\ else
                           \c$~<~Out_case_alt_30\;

  x2_64 <= resPtr_31;

  with (\c$~<~Out_case_scrut_63\(128 downto 128)) select
    \c$~<~Out_case_alt_30\ <= ( Tup2_sel0_signed => resPtr_31
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_32)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_31
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_32)
                               & std_logic_vector(x2_65 + to_signed(1,64))))) ) when others;

  x2_65 <= y_63;

  y_63 <= a1_30.Tup2_1_sel1_signed_1;

  a1_30 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_63\(127 downto 0)));

  -- index begin
  indexVec_63 : block
    signal vec_index_63 : integer range 0 to 64-1;
  begin
    vec_index_63 <= to_integer(resPtr_31)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_63\ <= currRes_31(vec_index_63);
  end block;
  -- index end

  currRes_31 <= \c$countConOut_app_arg_31\.Tup2_0_sel1_array_of_Maybe;

  resPtr_31 <= \c$countConOut_app_arg_31\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_64\ <= tagToEnum(\c$~<~Out_app_arg_65\);

  \c$~<~Out_app_arg_65\ <= to_signed(1,64) when x1_31 /= y_64 else to_signed(0,64);

  y_64 <= wild2_32;

  x1_31 <= wild2_31;

  -- index begin
  indexVec_64 : block
    signal vec_index_64 : integer range 0 to 64-1;
  begin
    vec_index_64 <= to_integer(to_signed(31,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_31 <= \c$app_arg\(vec_index_64);
  end block;
  -- index end

  \c$countConOut_app_arg_31\ <= ( Tup2_0_sel0_signed => x2_66 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_32\ ) when \c$~<~Out_case_scrut_66\ else
                                ( Tup2_0_sel0_signed => resPtr_32
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_32\ );

  clash_internal_cOut_32 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_32\
      , xs           => currRes_32
      , ds           => \c$~<~Out_app_arg_66\ );

  \c$~<~Out_app_arg_66\ <= ( Tup2_sel0_signed => x2_66 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_32)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_66\ else
                           \c$~<~Out_case_alt_31\;

  x2_66 <= resPtr_32;

  with (\c$~<~Out_case_scrut_65\(128 downto 128)) select
    \c$~<~Out_case_alt_31\ <= ( Tup2_sel0_signed => resPtr_32
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_33)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_32
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_33)
                               & std_logic_vector(x2_67 + to_signed(1,64))))) ) when others;

  x2_67 <= y_65;

  y_65 <= a1_31.Tup2_1_sel1_signed_1;

  a1_31 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_65\(127 downto 0)));

  -- index begin
  indexVec_65 : block
    signal vec_index_65 : integer range 0 to 64-1;
  begin
    vec_index_65 <= to_integer(resPtr_32)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_65\ <= currRes_32(vec_index_65);
  end block;
  -- index end

  currRes_32 <= \c$countConOut_app_arg_32\.Tup2_0_sel1_array_of_Maybe;

  resPtr_32 <= \c$countConOut_app_arg_32\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_66\ <= tagToEnum(\c$~<~Out_app_arg_67\);

  \c$~<~Out_app_arg_67\ <= to_signed(1,64) when x1_32 /= y_66 else to_signed(0,64);

  y_66 <= wild2_33;

  x1_32 <= wild2_32;

  -- index begin
  indexVec_66 : block
    signal vec_index_66 : integer range 0 to 64-1;
  begin
    vec_index_66 <= to_integer(to_signed(30,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_32 <= \c$app_arg\(vec_index_66);
  end block;
  -- index end

  \c$countConOut_app_arg_32\ <= ( Tup2_0_sel0_signed => x2_68 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_33\ ) when \c$~<~Out_case_scrut_68\ else
                                ( Tup2_0_sel0_signed => resPtr_33
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_33\ );

  clash_internal_cOut_33 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_33\
      , xs           => currRes_33
      , ds           => \c$~<~Out_app_arg_68\ );

  \c$~<~Out_app_arg_68\ <= ( Tup2_sel0_signed => x2_68 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_33)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_68\ else
                           \c$~<~Out_case_alt_32\;

  x2_68 <= resPtr_33;

  with (\c$~<~Out_case_scrut_67\(128 downto 128)) select
    \c$~<~Out_case_alt_32\ <= ( Tup2_sel0_signed => resPtr_33
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_34)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_33
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_34)
                               & std_logic_vector(x2_69 + to_signed(1,64))))) ) when others;

  x2_69 <= y_67;

  y_67 <= a1_32.Tup2_1_sel1_signed_1;

  a1_32 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_67\(127 downto 0)));

  -- index begin
  indexVec_67 : block
    signal vec_index_67 : integer range 0 to 64-1;
  begin
    vec_index_67 <= to_integer(resPtr_33)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_67\ <= currRes_33(vec_index_67);
  end block;
  -- index end

  currRes_33 <= \c$countConOut_app_arg_33\.Tup2_0_sel1_array_of_Maybe;

  resPtr_33 <= \c$countConOut_app_arg_33\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_68\ <= tagToEnum(\c$~<~Out_app_arg_69\);

  \c$~<~Out_app_arg_69\ <= to_signed(1,64) when x1_33 /= y_68 else to_signed(0,64);

  y_68 <= wild2_34;

  x1_33 <= wild2_33;

  -- index begin
  indexVec_68 : block
    signal vec_index_68 : integer range 0 to 64-1;
  begin
    vec_index_68 <= to_integer(to_signed(29,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_33 <= \c$app_arg\(vec_index_68);
  end block;
  -- index end

  \c$countConOut_app_arg_33\ <= ( Tup2_0_sel0_signed => x2_70 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_34\ ) when \c$~<~Out_case_scrut_70\ else
                                ( Tup2_0_sel0_signed => resPtr_34
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_34\ );

  clash_internal_cOut_34 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_34\
      , xs           => currRes_34
      , ds           => \c$~<~Out_app_arg_70\ );

  \c$~<~Out_app_arg_70\ <= ( Tup2_sel0_signed => x2_70 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_34)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_70\ else
                           \c$~<~Out_case_alt_33\;

  x2_70 <= resPtr_34;

  with (\c$~<~Out_case_scrut_69\(128 downto 128)) select
    \c$~<~Out_case_alt_33\ <= ( Tup2_sel0_signed => resPtr_34
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_35)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_34
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_35)
                               & std_logic_vector(x2_71 + to_signed(1,64))))) ) when others;

  x2_71 <= y_69;

  y_69 <= a1_33.Tup2_1_sel1_signed_1;

  a1_33 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_69\(127 downto 0)));

  -- index begin
  indexVec_69 : block
    signal vec_index_69 : integer range 0 to 64-1;
  begin
    vec_index_69 <= to_integer(resPtr_34)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_69\ <= currRes_34(vec_index_69);
  end block;
  -- index end

  currRes_34 <= \c$countConOut_app_arg_34\.Tup2_0_sel1_array_of_Maybe;

  resPtr_34 <= \c$countConOut_app_arg_34\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_70\ <= tagToEnum(\c$~<~Out_app_arg_71\);

  \c$~<~Out_app_arg_71\ <= to_signed(1,64) when x1_34 /= y_70 else to_signed(0,64);

  y_70 <= wild2_35;

  x1_34 <= wild2_34;

  -- index begin
  indexVec_70 : block
    signal vec_index_70 : integer range 0 to 64-1;
  begin
    vec_index_70 <= to_integer(to_signed(28,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_34 <= \c$app_arg\(vec_index_70);
  end block;
  -- index end

  \c$countConOut_app_arg_34\ <= ( Tup2_0_sel0_signed => x2_72 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_35\ ) when \c$~<~Out_case_scrut_72\ else
                                ( Tup2_0_sel0_signed => resPtr_35
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_35\ );

  clash_internal_cOut_35 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_35\
      , xs           => currRes_35
      , ds           => \c$~<~Out_app_arg_72\ );

  \c$~<~Out_app_arg_72\ <= ( Tup2_sel0_signed => x2_72 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_35)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_72\ else
                           \c$~<~Out_case_alt_34\;

  x2_72 <= resPtr_35;

  with (\c$~<~Out_case_scrut_71\(128 downto 128)) select
    \c$~<~Out_case_alt_34\ <= ( Tup2_sel0_signed => resPtr_35
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_36)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_35
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_36)
                               & std_logic_vector(x2_73 + to_signed(1,64))))) ) when others;

  x2_73 <= y_71;

  y_71 <= a1_34.Tup2_1_sel1_signed_1;

  a1_34 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_71\(127 downto 0)));

  -- index begin
  indexVec_71 : block
    signal vec_index_71 : integer range 0 to 64-1;
  begin
    vec_index_71 <= to_integer(resPtr_35)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_71\ <= currRes_35(vec_index_71);
  end block;
  -- index end

  currRes_35 <= \c$countConOut_app_arg_35\.Tup2_0_sel1_array_of_Maybe;

  resPtr_35 <= \c$countConOut_app_arg_35\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_72\ <= tagToEnum(\c$~<~Out_app_arg_73\);

  \c$~<~Out_app_arg_73\ <= to_signed(1,64) when x1_35 /= y_72 else to_signed(0,64);

  y_72 <= wild2_36;

  x1_35 <= wild2_35;

  -- index begin
  indexVec_72 : block
    signal vec_index_72 : integer range 0 to 64-1;
  begin
    vec_index_72 <= to_integer(to_signed(27,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_35 <= \c$app_arg\(vec_index_72);
  end block;
  -- index end

  \c$countConOut_app_arg_35\ <= ( Tup2_0_sel0_signed => x2_74 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_36\ ) when \c$~<~Out_case_scrut_74\ else
                                ( Tup2_0_sel0_signed => resPtr_36
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_36\ );

  clash_internal_cOut_36 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_36\
      , xs           => currRes_36
      , ds           => \c$~<~Out_app_arg_74\ );

  \c$~<~Out_app_arg_74\ <= ( Tup2_sel0_signed => x2_74 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_36)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_74\ else
                           \c$~<~Out_case_alt_35\;

  x2_74 <= resPtr_36;

  with (\c$~<~Out_case_scrut_73\(128 downto 128)) select
    \c$~<~Out_case_alt_35\ <= ( Tup2_sel0_signed => resPtr_36
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_37)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_36
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_37)
                               & std_logic_vector(x2_75 + to_signed(1,64))))) ) when others;

  x2_75 <= y_73;

  y_73 <= a1_35.Tup2_1_sel1_signed_1;

  a1_35 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_73\(127 downto 0)));

  -- index begin
  indexVec_73 : block
    signal vec_index_73 : integer range 0 to 64-1;
  begin
    vec_index_73 <= to_integer(resPtr_36)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_73\ <= currRes_36(vec_index_73);
  end block;
  -- index end

  currRes_36 <= \c$countConOut_app_arg_36\.Tup2_0_sel1_array_of_Maybe;

  resPtr_36 <= \c$countConOut_app_arg_36\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_74\ <= tagToEnum(\c$~<~Out_app_arg_75\);

  \c$~<~Out_app_arg_75\ <= to_signed(1,64) when x1_36 /= y_74 else to_signed(0,64);

  y_74 <= wild2_37;

  x1_36 <= wild2_36;

  -- index begin
  indexVec_74 : block
    signal vec_index_74 : integer range 0 to 64-1;
  begin
    vec_index_74 <= to_integer(to_signed(26,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_36 <= \c$app_arg\(vec_index_74);
  end block;
  -- index end

  \c$countConOut_app_arg_36\ <= ( Tup2_0_sel0_signed => x2_76 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_37\ ) when \c$~<~Out_case_scrut_76\ else
                                ( Tup2_0_sel0_signed => resPtr_37
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_37\ );

  clash_internal_cOut_37 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_37\
      , xs           => currRes_37
      , ds           => \c$~<~Out_app_arg_76\ );

  \c$~<~Out_app_arg_76\ <= ( Tup2_sel0_signed => x2_76 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_37)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_76\ else
                           \c$~<~Out_case_alt_36\;

  x2_76 <= resPtr_37;

  with (\c$~<~Out_case_scrut_75\(128 downto 128)) select
    \c$~<~Out_case_alt_36\ <= ( Tup2_sel0_signed => resPtr_37
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_38)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_37
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_38)
                               & std_logic_vector(x2_77 + to_signed(1,64))))) ) when others;

  x2_77 <= y_75;

  y_75 <= a1_36.Tup2_1_sel1_signed_1;

  a1_36 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_75\(127 downto 0)));

  -- index begin
  indexVec_75 : block
    signal vec_index_75 : integer range 0 to 64-1;
  begin
    vec_index_75 <= to_integer(resPtr_37)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_75\ <= currRes_37(vec_index_75);
  end block;
  -- index end

  currRes_37 <= \c$countConOut_app_arg_37\.Tup2_0_sel1_array_of_Maybe;

  resPtr_37 <= \c$countConOut_app_arg_37\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_76\ <= tagToEnum(\c$~<~Out_app_arg_77\);

  \c$~<~Out_app_arg_77\ <= to_signed(1,64) when x1_37 /= y_76 else to_signed(0,64);

  y_76 <= wild2_38;

  x1_37 <= wild2_37;

  -- index begin
  indexVec_76 : block
    signal vec_index_76 : integer range 0 to 64-1;
  begin
    vec_index_76 <= to_integer(to_signed(25,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_37 <= \c$app_arg\(vec_index_76);
  end block;
  -- index end

  \c$countConOut_app_arg_37\ <= ( Tup2_0_sel0_signed => x2_78 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_38\ ) when \c$~<~Out_case_scrut_78\ else
                                ( Tup2_0_sel0_signed => resPtr_38
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_38\ );

  clash_internal_cOut_38 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_38\
      , xs           => currRes_38
      , ds           => \c$~<~Out_app_arg_78\ );

  \c$~<~Out_app_arg_78\ <= ( Tup2_sel0_signed => x2_78 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_38)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_78\ else
                           \c$~<~Out_case_alt_37\;

  x2_78 <= resPtr_38;

  with (\c$~<~Out_case_scrut_77\(128 downto 128)) select
    \c$~<~Out_case_alt_37\ <= ( Tup2_sel0_signed => resPtr_38
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_39)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_38
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_39)
                               & std_logic_vector(x2_79 + to_signed(1,64))))) ) when others;

  x2_79 <= y_77;

  y_77 <= a1_37.Tup2_1_sel1_signed_1;

  a1_37 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_77\(127 downto 0)));

  -- index begin
  indexVec_77 : block
    signal vec_index_77 : integer range 0 to 64-1;
  begin
    vec_index_77 <= to_integer(resPtr_38)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_77\ <= currRes_38(vec_index_77);
  end block;
  -- index end

  currRes_38 <= \c$countConOut_app_arg_38\.Tup2_0_sel1_array_of_Maybe;

  resPtr_38 <= \c$countConOut_app_arg_38\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_78\ <= tagToEnum(\c$~<~Out_app_arg_79\);

  \c$~<~Out_app_arg_79\ <= to_signed(1,64) when x1_38 /= y_78 else to_signed(0,64);

  y_78 <= wild2_39;

  x1_38 <= wild2_38;

  -- index begin
  indexVec_78 : block
    signal vec_index_78 : integer range 0 to 64-1;
  begin
    vec_index_78 <= to_integer(to_signed(24,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_38 <= \c$app_arg\(vec_index_78);
  end block;
  -- index end

  \c$countConOut_app_arg_38\ <= ( Tup2_0_sel0_signed => x2_80 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_39\ ) when \c$~<~Out_case_scrut_80\ else
                                ( Tup2_0_sel0_signed => resPtr_39
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_39\ );

  clash_internal_cOut_39 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_39\
      , xs           => currRes_39
      , ds           => \c$~<~Out_app_arg_80\ );

  \c$~<~Out_app_arg_80\ <= ( Tup2_sel0_signed => x2_80 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_39)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_80\ else
                           \c$~<~Out_case_alt_38\;

  x2_80 <= resPtr_39;

  with (\c$~<~Out_case_scrut_79\(128 downto 128)) select
    \c$~<~Out_case_alt_38\ <= ( Tup2_sel0_signed => resPtr_39
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_40)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_39
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_40)
                               & std_logic_vector(x2_81 + to_signed(1,64))))) ) when others;

  x2_81 <= y_79;

  y_79 <= a1_38.Tup2_1_sel1_signed_1;

  a1_38 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_79\(127 downto 0)));

  -- index begin
  indexVec_79 : block
    signal vec_index_79 : integer range 0 to 64-1;
  begin
    vec_index_79 <= to_integer(resPtr_39)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_79\ <= currRes_39(vec_index_79);
  end block;
  -- index end

  currRes_39 <= \c$countConOut_app_arg_39\.Tup2_0_sel1_array_of_Maybe;

  resPtr_39 <= \c$countConOut_app_arg_39\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_80\ <= tagToEnum(\c$~<~Out_app_arg_81\);

  \c$~<~Out_app_arg_81\ <= to_signed(1,64) when x1_39 /= y_80 else to_signed(0,64);

  y_80 <= wild2_40;

  x1_39 <= wild2_39;

  -- index begin
  indexVec_80 : block
    signal vec_index_80 : integer range 0 to 64-1;
  begin
    vec_index_80 <= to_integer(to_signed(23,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_39 <= \c$app_arg\(vec_index_80);
  end block;
  -- index end

  \c$countConOut_app_arg_39\ <= ( Tup2_0_sel0_signed => x2_82 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_40\ ) when \c$~<~Out_case_scrut_82\ else
                                ( Tup2_0_sel0_signed => resPtr_40
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_40\ );

  clash_internal_cOut_40 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_40\
      , xs           => currRes_40
      , ds           => \c$~<~Out_app_arg_82\ );

  \c$~<~Out_app_arg_82\ <= ( Tup2_sel0_signed => x2_82 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_40)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_82\ else
                           \c$~<~Out_case_alt_39\;

  x2_82 <= resPtr_40;

  with (\c$~<~Out_case_scrut_81\(128 downto 128)) select
    \c$~<~Out_case_alt_39\ <= ( Tup2_sel0_signed => resPtr_40
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_41)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_40
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_41)
                               & std_logic_vector(x2_83 + to_signed(1,64))))) ) when others;

  x2_83 <= y_81;

  y_81 <= a1_39.Tup2_1_sel1_signed_1;

  a1_39 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_81\(127 downto 0)));

  -- index begin
  indexVec_81 : block
    signal vec_index_81 : integer range 0 to 64-1;
  begin
    vec_index_81 <= to_integer(resPtr_40)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_81\ <= currRes_40(vec_index_81);
  end block;
  -- index end

  currRes_40 <= \c$countConOut_app_arg_40\.Tup2_0_sel1_array_of_Maybe;

  resPtr_40 <= \c$countConOut_app_arg_40\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_82\ <= tagToEnum(\c$~<~Out_app_arg_83\);

  \c$~<~Out_app_arg_83\ <= to_signed(1,64) when x1_40 /= y_82 else to_signed(0,64);

  y_82 <= wild2_41;

  x1_40 <= wild2_40;

  -- index begin
  indexVec_82 : block
    signal vec_index_82 : integer range 0 to 64-1;
  begin
    vec_index_82 <= to_integer(to_signed(22,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_40 <= \c$app_arg\(vec_index_82);
  end block;
  -- index end

  \c$countConOut_app_arg_40\ <= ( Tup2_0_sel0_signed => x2_84 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_41\ ) when \c$~<~Out_case_scrut_84\ else
                                ( Tup2_0_sel0_signed => resPtr_41
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_41\ );

  clash_internal_cOut_41 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_41\
      , xs           => currRes_41
      , ds           => \c$~<~Out_app_arg_84\ );

  \c$~<~Out_app_arg_84\ <= ( Tup2_sel0_signed => x2_84 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_41)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_84\ else
                           \c$~<~Out_case_alt_40\;

  x2_84 <= resPtr_41;

  with (\c$~<~Out_case_scrut_83\(128 downto 128)) select
    \c$~<~Out_case_alt_40\ <= ( Tup2_sel0_signed => resPtr_41
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_42)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_41
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_42)
                               & std_logic_vector(x2_85 + to_signed(1,64))))) ) when others;

  x2_85 <= y_83;

  y_83 <= a1_40.Tup2_1_sel1_signed_1;

  a1_40 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_83\(127 downto 0)));

  -- index begin
  indexVec_83 : block
    signal vec_index_83 : integer range 0 to 64-1;
  begin
    vec_index_83 <= to_integer(resPtr_41)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_83\ <= currRes_41(vec_index_83);
  end block;
  -- index end

  currRes_41 <= \c$countConOut_app_arg_41\.Tup2_0_sel1_array_of_Maybe;

  resPtr_41 <= \c$countConOut_app_arg_41\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_84\ <= tagToEnum(\c$~<~Out_app_arg_85\);

  \c$~<~Out_app_arg_85\ <= to_signed(1,64) when x1_41 /= y_84 else to_signed(0,64);

  y_84 <= wild2_42;

  x1_41 <= wild2_41;

  -- index begin
  indexVec_84 : block
    signal vec_index_84 : integer range 0 to 64-1;
  begin
    vec_index_84 <= to_integer(to_signed(21,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_41 <= \c$app_arg\(vec_index_84);
  end block;
  -- index end

  \c$countConOut_app_arg_41\ <= ( Tup2_0_sel0_signed => x2_86 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_42\ ) when \c$~<~Out_case_scrut_86\ else
                                ( Tup2_0_sel0_signed => resPtr_42
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_42\ );

  clash_internal_cOut_42 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_42\
      , xs           => currRes_42
      , ds           => \c$~<~Out_app_arg_86\ );

  \c$~<~Out_app_arg_86\ <= ( Tup2_sel0_signed => x2_86 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_42)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_86\ else
                           \c$~<~Out_case_alt_41\;

  x2_86 <= resPtr_42;

  with (\c$~<~Out_case_scrut_85\(128 downto 128)) select
    \c$~<~Out_case_alt_41\ <= ( Tup2_sel0_signed => resPtr_42
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_43)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_42
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_43)
                               & std_logic_vector(x2_87 + to_signed(1,64))))) ) when others;

  x2_87 <= y_85;

  y_85 <= a1_41.Tup2_1_sel1_signed_1;

  a1_41 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_85\(127 downto 0)));

  -- index begin
  indexVec_85 : block
    signal vec_index_85 : integer range 0 to 64-1;
  begin
    vec_index_85 <= to_integer(resPtr_42)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_85\ <= currRes_42(vec_index_85);
  end block;
  -- index end

  currRes_42 <= \c$countConOut_app_arg_42\.Tup2_0_sel1_array_of_Maybe;

  resPtr_42 <= \c$countConOut_app_arg_42\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_86\ <= tagToEnum(\c$~<~Out_app_arg_87\);

  \c$~<~Out_app_arg_87\ <= to_signed(1,64) when x1_42 /= y_86 else to_signed(0,64);

  y_86 <= wild2_43;

  x1_42 <= wild2_42;

  -- index begin
  indexVec_86 : block
    signal vec_index_86 : integer range 0 to 64-1;
  begin
    vec_index_86 <= to_integer(to_signed(20,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_42 <= \c$app_arg\(vec_index_86);
  end block;
  -- index end

  \c$countConOut_app_arg_42\ <= ( Tup2_0_sel0_signed => x2_88 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_43\ ) when \c$~<~Out_case_scrut_88\ else
                                ( Tup2_0_sel0_signed => resPtr_43
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_43\ );

  clash_internal_cOut_43 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_43\
      , xs           => currRes_43
      , ds           => \c$~<~Out_app_arg_88\ );

  \c$~<~Out_app_arg_88\ <= ( Tup2_sel0_signed => x2_88 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_43)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_88\ else
                           \c$~<~Out_case_alt_42\;

  x2_88 <= resPtr_43;

  with (\c$~<~Out_case_scrut_87\(128 downto 128)) select
    \c$~<~Out_case_alt_42\ <= ( Tup2_sel0_signed => resPtr_43
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_44)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_43
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_44)
                               & std_logic_vector(x2_89 + to_signed(1,64))))) ) when others;

  x2_89 <= y_87;

  y_87 <= a1_42.Tup2_1_sel1_signed_1;

  a1_42 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_87\(127 downto 0)));

  -- index begin
  indexVec_87 : block
    signal vec_index_87 : integer range 0 to 64-1;
  begin
    vec_index_87 <= to_integer(resPtr_43)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_87\ <= currRes_43(vec_index_87);
  end block;
  -- index end

  currRes_43 <= \c$countConOut_app_arg_43\.Tup2_0_sel1_array_of_Maybe;

  resPtr_43 <= \c$countConOut_app_arg_43\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_88\ <= tagToEnum(\c$~<~Out_app_arg_89\);

  \c$~<~Out_app_arg_89\ <= to_signed(1,64) when x1_43 /= y_88 else to_signed(0,64);

  y_88 <= wild2_44;

  x1_43 <= wild2_43;

  -- index begin
  indexVec_88 : block
    signal vec_index_88 : integer range 0 to 64-1;
  begin
    vec_index_88 <= to_integer(to_signed(19,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_43 <= \c$app_arg\(vec_index_88);
  end block;
  -- index end

  \c$countConOut_app_arg_43\ <= ( Tup2_0_sel0_signed => x2_90 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_44\ ) when \c$~<~Out_case_scrut_90\ else
                                ( Tup2_0_sel0_signed => resPtr_44
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_44\ );

  clash_internal_cOut_44 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_44\
      , xs           => currRes_44
      , ds           => \c$~<~Out_app_arg_90\ );

  \c$~<~Out_app_arg_90\ <= ( Tup2_sel0_signed => x2_90 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_44)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_90\ else
                           \c$~<~Out_case_alt_43\;

  x2_90 <= resPtr_44;

  with (\c$~<~Out_case_scrut_89\(128 downto 128)) select
    \c$~<~Out_case_alt_43\ <= ( Tup2_sel0_signed => resPtr_44
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_45)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_44
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_45)
                               & std_logic_vector(x2_91 + to_signed(1,64))))) ) when others;

  x2_91 <= y_89;

  y_89 <= a1_43.Tup2_1_sel1_signed_1;

  a1_43 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_89\(127 downto 0)));

  -- index begin
  indexVec_89 : block
    signal vec_index_89 : integer range 0 to 64-1;
  begin
    vec_index_89 <= to_integer(resPtr_44)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_89\ <= currRes_44(vec_index_89);
  end block;
  -- index end

  currRes_44 <= \c$countConOut_app_arg_44\.Tup2_0_sel1_array_of_Maybe;

  resPtr_44 <= \c$countConOut_app_arg_44\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_90\ <= tagToEnum(\c$~<~Out_app_arg_91\);

  \c$~<~Out_app_arg_91\ <= to_signed(1,64) when x1_44 /= y_90 else to_signed(0,64);

  y_90 <= wild2_45;

  x1_44 <= wild2_44;

  -- index begin
  indexVec_90 : block
    signal vec_index_90 : integer range 0 to 64-1;
  begin
    vec_index_90 <= to_integer(to_signed(18,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_44 <= \c$app_arg\(vec_index_90);
  end block;
  -- index end

  \c$countConOut_app_arg_44\ <= ( Tup2_0_sel0_signed => x2_92 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_45\ ) when \c$~<~Out_case_scrut_92\ else
                                ( Tup2_0_sel0_signed => resPtr_45
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_45\ );

  clash_internal_cOut_45 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_45\
      , xs           => currRes_45
      , ds           => \c$~<~Out_app_arg_92\ );

  \c$~<~Out_app_arg_92\ <= ( Tup2_sel0_signed => x2_92 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_45)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_92\ else
                           \c$~<~Out_case_alt_44\;

  x2_92 <= resPtr_45;

  with (\c$~<~Out_case_scrut_91\(128 downto 128)) select
    \c$~<~Out_case_alt_44\ <= ( Tup2_sel0_signed => resPtr_45
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_46)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_45
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_46)
                               & std_logic_vector(x2_93 + to_signed(1,64))))) ) when others;

  x2_93 <= y_91;

  y_91 <= a1_44.Tup2_1_sel1_signed_1;

  a1_44 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_91\(127 downto 0)));

  -- index begin
  indexVec_91 : block
    signal vec_index_91 : integer range 0 to 64-1;
  begin
    vec_index_91 <= to_integer(resPtr_45)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_91\ <= currRes_45(vec_index_91);
  end block;
  -- index end

  currRes_45 <= \c$countConOut_app_arg_45\.Tup2_0_sel1_array_of_Maybe;

  resPtr_45 <= \c$countConOut_app_arg_45\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_92\ <= tagToEnum(\c$~<~Out_app_arg_93\);

  \c$~<~Out_app_arg_93\ <= to_signed(1,64) when x1_45 /= y_92 else to_signed(0,64);

  y_92 <= wild2_46;

  x1_45 <= wild2_45;

  -- index begin
  indexVec_92 : block
    signal vec_index_92 : integer range 0 to 64-1;
  begin
    vec_index_92 <= to_integer(to_signed(17,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_45 <= \c$app_arg\(vec_index_92);
  end block;
  -- index end

  \c$countConOut_app_arg_45\ <= ( Tup2_0_sel0_signed => x2_94 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_46\ ) when \c$~<~Out_case_scrut_94\ else
                                ( Tup2_0_sel0_signed => resPtr_46
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_46\ );

  clash_internal_cOut_46 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_46\
      , xs           => currRes_46
      , ds           => \c$~<~Out_app_arg_94\ );

  \c$~<~Out_app_arg_94\ <= ( Tup2_sel0_signed => x2_94 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_46)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_94\ else
                           \c$~<~Out_case_alt_45\;

  x2_94 <= resPtr_46;

  with (\c$~<~Out_case_scrut_93\(128 downto 128)) select
    \c$~<~Out_case_alt_45\ <= ( Tup2_sel0_signed => resPtr_46
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_47)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_46
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_47)
                               & std_logic_vector(x2_95 + to_signed(1,64))))) ) when others;

  x2_95 <= y_93;

  y_93 <= a1_45.Tup2_1_sel1_signed_1;

  a1_45 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_93\(127 downto 0)));

  -- index begin
  indexVec_93 : block
    signal vec_index_93 : integer range 0 to 64-1;
  begin
    vec_index_93 <= to_integer(resPtr_46)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_93\ <= currRes_46(vec_index_93);
  end block;
  -- index end

  currRes_46 <= \c$countConOut_app_arg_46\.Tup2_0_sel1_array_of_Maybe;

  resPtr_46 <= \c$countConOut_app_arg_46\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_94\ <= tagToEnum(\c$~<~Out_app_arg_95\);

  \c$~<~Out_app_arg_95\ <= to_signed(1,64) when x1_46 /= y_94 else to_signed(0,64);

  y_94 <= wild2_47;

  x1_46 <= wild2_46;

  -- index begin
  indexVec_94 : block
    signal vec_index_94 : integer range 0 to 64-1;
  begin
    vec_index_94 <= to_integer(to_signed(16,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_46 <= \c$app_arg\(vec_index_94);
  end block;
  -- index end

  \c$countConOut_app_arg_46\ <= ( Tup2_0_sel0_signed => x2_96 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_47\ ) when \c$~<~Out_case_scrut_96\ else
                                ( Tup2_0_sel0_signed => resPtr_47
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_47\ );

  clash_internal_cOut_47 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_47\
      , xs           => currRes_47
      , ds           => \c$~<~Out_app_arg_96\ );

  \c$~<~Out_app_arg_96\ <= ( Tup2_sel0_signed => x2_96 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_47)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_96\ else
                           \c$~<~Out_case_alt_46\;

  x2_96 <= resPtr_47;

  with (\c$~<~Out_case_scrut_95\(128 downto 128)) select
    \c$~<~Out_case_alt_46\ <= ( Tup2_sel0_signed => resPtr_47
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_48)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_47
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_48)
                               & std_logic_vector(x2_97 + to_signed(1,64))))) ) when others;

  x2_97 <= y_95;

  y_95 <= a1_46.Tup2_1_sel1_signed_1;

  a1_46 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_95\(127 downto 0)));

  -- index begin
  indexVec_95 : block
    signal vec_index_95 : integer range 0 to 64-1;
  begin
    vec_index_95 <= to_integer(resPtr_47)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_95\ <= currRes_47(vec_index_95);
  end block;
  -- index end

  currRes_47 <= \c$countConOut_app_arg_47\.Tup2_0_sel1_array_of_Maybe;

  resPtr_47 <= \c$countConOut_app_arg_47\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_96\ <= tagToEnum(\c$~<~Out_app_arg_97\);

  \c$~<~Out_app_arg_97\ <= to_signed(1,64) when x1_47 /= y_96 else to_signed(0,64);

  y_96 <= wild2_48;

  x1_47 <= wild2_47;

  -- index begin
  indexVec_96 : block
    signal vec_index_96 : integer range 0 to 64-1;
  begin
    vec_index_96 <= to_integer(to_signed(15,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_47 <= \c$app_arg\(vec_index_96);
  end block;
  -- index end

  \c$countConOut_app_arg_47\ <= ( Tup2_0_sel0_signed => x2_98 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_48\ ) when \c$~<~Out_case_scrut_98\ else
                                ( Tup2_0_sel0_signed => resPtr_48
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_48\ );

  clash_internal_cOut_48 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_48\
      , xs           => currRes_48
      , ds           => \c$~<~Out_app_arg_98\ );

  \c$~<~Out_app_arg_98\ <= ( Tup2_sel0_signed => x2_98 + to_signed(1,64)
                           , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_48)
                            & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_98\ else
                           \c$~<~Out_case_alt_47\;

  x2_98 <= resPtr_48;

  with (\c$~<~Out_case_scrut_97\(128 downto 128)) select
    \c$~<~Out_case_alt_47\ <= ( Tup2_sel0_signed => resPtr_48
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_49)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_48
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_49)
                               & std_logic_vector(x2_99 + to_signed(1,64))))) ) when others;

  x2_99 <= y_97;

  y_97 <= a1_47.Tup2_1_sel1_signed_1;

  a1_47 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_97\(127 downto 0)));

  -- index begin
  indexVec_97 : block
    signal vec_index_97 : integer range 0 to 64-1;
  begin
    vec_index_97 <= to_integer(resPtr_48)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_97\ <= currRes_48(vec_index_97);
  end block;
  -- index end

  currRes_48 <= \c$countConOut_app_arg_48\.Tup2_0_sel1_array_of_Maybe;

  resPtr_48 <= \c$countConOut_app_arg_48\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_98\ <= tagToEnum(\c$~<~Out_app_arg_99\);

  \c$~<~Out_app_arg_99\ <= to_signed(1,64) when x1_48 /= y_98 else to_signed(0,64);

  y_98 <= wild2_49;

  x1_48 <= wild2_48;

  -- index begin
  indexVec_98 : block
    signal vec_index_98 : integer range 0 to 64-1;
  begin
    vec_index_98 <= to_integer(to_signed(14,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_48 <= \c$app_arg\(vec_index_98);
  end block;
  -- index end

  \c$countConOut_app_arg_48\ <= ( Tup2_0_sel0_signed => x2_100 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_49\ ) when \c$~<~Out_case_scrut_100\ else
                                ( Tup2_0_sel0_signed => resPtr_49
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_49\ );

  clash_internal_cOut_49 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_49\
      , xs           => currRes_49
      , ds           => \c$~<~Out_app_arg_100\ );

  \c$~<~Out_app_arg_100\ <= ( Tup2_sel0_signed => x2_100 + to_signed(1,64)
                            , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_49)
                             & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_100\ else
                            \c$~<~Out_case_alt_48\;

  x2_100 <= resPtr_49;

  with (\c$~<~Out_case_scrut_99\(128 downto 128)) select
    \c$~<~Out_case_alt_48\ <= ( Tup2_sel0_signed => resPtr_49
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_50)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_49
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_50)
                               & std_logic_vector(x2_101 + to_signed(1,64))))) ) when others;

  x2_101 <= y_99;

  y_99 <= a1_48.Tup2_1_sel1_signed_1;

  a1_48 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_99\(127 downto 0)));

  -- index begin
  indexVec_99 : block
    signal vec_index_99 : integer range 0 to 64-1;
  begin
    vec_index_99 <= to_integer(resPtr_49)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_99\ <= currRes_49(vec_index_99);
  end block;
  -- index end

  currRes_49 <= \c$countConOut_app_arg_49\.Tup2_0_sel1_array_of_Maybe;

  resPtr_49 <= \c$countConOut_app_arg_49\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_100\ <= tagToEnum(\c$~<~Out_app_arg_101\);

  \c$~<~Out_app_arg_101\ <= to_signed(1,64) when x1_49 /= y_100 else to_signed(0,64);

  y_100 <= wild2_50;

  x1_49 <= wild2_49;

  -- index begin
  indexVec_100 : block
    signal vec_index_100 : integer range 0 to 64-1;
  begin
    vec_index_100 <= to_integer(to_signed(13,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_49 <= \c$app_arg\(vec_index_100);
  end block;
  -- index end

  \c$countConOut_app_arg_49\ <= ( Tup2_0_sel0_signed => x2_102 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_50\ ) when \c$~<~Out_case_scrut_102\ else
                                ( Tup2_0_sel0_signed => resPtr_50
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_50\ );

  clash_internal_cOut_50 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_50\
      , xs           => currRes_50
      , ds           => \c$~<~Out_app_arg_102\ );

  \c$~<~Out_app_arg_102\ <= ( Tup2_sel0_signed => x2_102 + to_signed(1,64)
                            , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_50)
                             & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_102\ else
                            \c$~<~Out_case_alt_49\;

  x2_102 <= resPtr_50;

  with (\c$~<~Out_case_scrut_101\(128 downto 128)) select
    \c$~<~Out_case_alt_49\ <= ( Tup2_sel0_signed => resPtr_50
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_51)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_50
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_51)
                               & std_logic_vector(x2_103 + to_signed(1,64))))) ) when others;

  x2_103 <= y_101;

  y_101 <= a1_49.Tup2_1_sel1_signed_1;

  a1_49 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_101\(127 downto 0)));

  -- index begin
  indexVec_101 : block
    signal vec_index_101 : integer range 0 to 64-1;
  begin
    vec_index_101 <= to_integer(resPtr_50)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_101\ <= currRes_50(vec_index_101);
  end block;
  -- index end

  currRes_50 <= \c$countConOut_app_arg_50\.Tup2_0_sel1_array_of_Maybe;

  resPtr_50 <= \c$countConOut_app_arg_50\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_102\ <= tagToEnum(\c$~<~Out_app_arg_103\);

  \c$~<~Out_app_arg_103\ <= to_signed(1,64) when x1_50 /= y_102 else to_signed(0,64);

  y_102 <= wild2_51;

  x1_50 <= wild2_50;

  -- index begin
  indexVec_102 : block
    signal vec_index_102 : integer range 0 to 64-1;
  begin
    vec_index_102 <= to_integer(to_signed(12,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_50 <= \c$app_arg\(vec_index_102);
  end block;
  -- index end

  \c$countConOut_app_arg_50\ <= ( Tup2_0_sel0_signed => x2_104 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_51\ ) when \c$~<~Out_case_scrut_104\ else
                                ( Tup2_0_sel0_signed => resPtr_51
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_51\ );

  clash_internal_cOut_51 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_51\
      , xs           => currRes_51
      , ds           => \c$~<~Out_app_arg_104\ );

  \c$~<~Out_app_arg_104\ <= ( Tup2_sel0_signed => x2_104 + to_signed(1,64)
                            , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_51)
                             & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_104\ else
                            \c$~<~Out_case_alt_50\;

  x2_104 <= resPtr_51;

  with (\c$~<~Out_case_scrut_103\(128 downto 128)) select
    \c$~<~Out_case_alt_50\ <= ( Tup2_sel0_signed => resPtr_51
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_52)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_51
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_52)
                               & std_logic_vector(x2_105 + to_signed(1,64))))) ) when others;

  x2_105 <= y_103;

  y_103 <= a1_50.Tup2_1_sel1_signed_1;

  a1_50 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_103\(127 downto 0)));

  -- index begin
  indexVec_103 : block
    signal vec_index_103 : integer range 0 to 64-1;
  begin
    vec_index_103 <= to_integer(resPtr_51)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_103\ <= currRes_51(vec_index_103);
  end block;
  -- index end

  currRes_51 <= \c$countConOut_app_arg_51\.Tup2_0_sel1_array_of_Maybe;

  resPtr_51 <= \c$countConOut_app_arg_51\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_104\ <= tagToEnum(\c$~<~Out_app_arg_105\);

  \c$~<~Out_app_arg_105\ <= to_signed(1,64) when x1_51 /= y_104 else to_signed(0,64);

  y_104 <= wild2_52;

  x1_51 <= wild2_51;

  -- index begin
  indexVec_104 : block
    signal vec_index_104 : integer range 0 to 64-1;
  begin
    vec_index_104 <= to_integer(to_signed(11,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_51 <= \c$app_arg\(vec_index_104);
  end block;
  -- index end

  \c$countConOut_app_arg_51\ <= ( Tup2_0_sel0_signed => x2_106 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_52\ ) when \c$~<~Out_case_scrut_106\ else
                                ( Tup2_0_sel0_signed => resPtr_52
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_52\ );

  clash_internal_cOut_52 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_52\
      , xs           => currRes_52
      , ds           => \c$~<~Out_app_arg_106\ );

  \c$~<~Out_app_arg_106\ <= ( Tup2_sel0_signed => x2_106 + to_signed(1,64)
                            , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_52)
                             & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_106\ else
                            \c$~<~Out_case_alt_51\;

  x2_106 <= resPtr_52;

  with (\c$~<~Out_case_scrut_105\(128 downto 128)) select
    \c$~<~Out_case_alt_51\ <= ( Tup2_sel0_signed => resPtr_52
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_53)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_52
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_53)
                               & std_logic_vector(x2_107 + to_signed(1,64))))) ) when others;

  x2_107 <= y_105;

  y_105 <= a1_51.Tup2_1_sel1_signed_1;

  a1_51 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_105\(127 downto 0)));

  -- index begin
  indexVec_105 : block
    signal vec_index_105 : integer range 0 to 64-1;
  begin
    vec_index_105 <= to_integer(resPtr_52)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_105\ <= currRes_52(vec_index_105);
  end block;
  -- index end

  currRes_52 <= \c$countConOut_app_arg_52\.Tup2_0_sel1_array_of_Maybe;

  resPtr_52 <= \c$countConOut_app_arg_52\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_106\ <= tagToEnum(\c$~<~Out_app_arg_107\);

  \c$~<~Out_app_arg_107\ <= to_signed(1,64) when x1_52 /= y_106 else to_signed(0,64);

  y_106 <= wild2_53;

  x1_52 <= wild2_52;

  -- index begin
  indexVec_106 : block
    signal vec_index_106 : integer range 0 to 64-1;
  begin
    vec_index_106 <= to_integer(to_signed(10,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_52 <= \c$app_arg\(vec_index_106);
  end block;
  -- index end

  \c$countConOut_app_arg_52\ <= ( Tup2_0_sel0_signed => x2_108 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_53\ ) when \c$~<~Out_case_scrut_108\ else
                                ( Tup2_0_sel0_signed => resPtr_53
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_53\ );

  clash_internal_cOut_53 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_53\
      , xs           => currRes_53
      , ds           => \c$~<~Out_app_arg_108\ );

  \c$~<~Out_app_arg_108\ <= ( Tup2_sel0_signed => x2_108 + to_signed(1,64)
                            , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_53)
                             & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_108\ else
                            \c$~<~Out_case_alt_52\;

  x2_108 <= resPtr_53;

  with (\c$~<~Out_case_scrut_107\(128 downto 128)) select
    \c$~<~Out_case_alt_52\ <= ( Tup2_sel0_signed => resPtr_53
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_54)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_53
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_54)
                               & std_logic_vector(x2_109 + to_signed(1,64))))) ) when others;

  x2_109 <= y_107;

  y_107 <= a1_52.Tup2_1_sel1_signed_1;

  a1_52 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_107\(127 downto 0)));

  -- index begin
  indexVec_107 : block
    signal vec_index_107 : integer range 0 to 64-1;
  begin
    vec_index_107 <= to_integer(resPtr_53)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_107\ <= currRes_53(vec_index_107);
  end block;
  -- index end

  currRes_53 <= \c$countConOut_app_arg_53\.Tup2_0_sel1_array_of_Maybe;

  resPtr_53 <= \c$countConOut_app_arg_53\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_108\ <= tagToEnum(\c$~<~Out_app_arg_109\);

  \c$~<~Out_app_arg_109\ <= to_signed(1,64) when x1_53 /= y_108 else to_signed(0,64);

  y_108 <= wild2_54;

  x1_53 <= wild2_53;

  -- index begin
  indexVec_108 : block
    signal vec_index_108 : integer range 0 to 64-1;
  begin
    vec_index_108 <= to_integer(to_signed(9,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_53 <= \c$app_arg\(vec_index_108);
  end block;
  -- index end

  \c$countConOut_app_arg_53\ <= ( Tup2_0_sel0_signed => x2_110 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_54\ ) when \c$~<~Out_case_scrut_110\ else
                                ( Tup2_0_sel0_signed => resPtr_54
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_54\ );

  clash_internal_cOut_54 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_54\
      , xs           => currRes_54
      , ds           => \c$~<~Out_app_arg_110\ );

  \c$~<~Out_app_arg_110\ <= ( Tup2_sel0_signed => x2_110 + to_signed(1,64)
                            , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_54)
                             & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_110\ else
                            \c$~<~Out_case_alt_53\;

  x2_110 <= resPtr_54;

  with (\c$~<~Out_case_scrut_109\(128 downto 128)) select
    \c$~<~Out_case_alt_53\ <= ( Tup2_sel0_signed => resPtr_54
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_55)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_54
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_55)
                               & std_logic_vector(x2_111 + to_signed(1,64))))) ) when others;

  x2_111 <= y_109;

  y_109 <= a1_53.Tup2_1_sel1_signed_1;

  a1_53 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_109\(127 downto 0)));

  -- index begin
  indexVec_109 : block
    signal vec_index_109 : integer range 0 to 64-1;
  begin
    vec_index_109 <= to_integer(resPtr_54)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_109\ <= currRes_54(vec_index_109);
  end block;
  -- index end

  currRes_54 <= \c$countConOut_app_arg_54\.Tup2_0_sel1_array_of_Maybe;

  resPtr_54 <= \c$countConOut_app_arg_54\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_110\ <= tagToEnum(\c$~<~Out_app_arg_111\);

  \c$~<~Out_app_arg_111\ <= to_signed(1,64) when x1_54 /= y_110 else to_signed(0,64);

  y_110 <= wild2_55;

  x1_54 <= wild2_54;

  -- index begin
  indexVec_110 : block
    signal vec_index_110 : integer range 0 to 64-1;
  begin
    vec_index_110 <= to_integer(to_signed(8,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_54 <= \c$app_arg\(vec_index_110);
  end block;
  -- index end

  \c$countConOut_app_arg_54\ <= ( Tup2_0_sel0_signed => x2_112 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_55\ ) when \c$~<~Out_case_scrut_112\ else
                                ( Tup2_0_sel0_signed => resPtr_55
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_55\ );

  clash_internal_cOut_55 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_55\
      , xs           => currRes_55
      , ds           => \c$~<~Out_app_arg_112\ );

  \c$~<~Out_app_arg_112\ <= ( Tup2_sel0_signed => x2_112 + to_signed(1,64)
                            , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_55)
                             & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_112\ else
                            \c$~<~Out_case_alt_54\;

  x2_112 <= resPtr_55;

  with (\c$~<~Out_case_scrut_111\(128 downto 128)) select
    \c$~<~Out_case_alt_54\ <= ( Tup2_sel0_signed => resPtr_55
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_56)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_55
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_56)
                               & std_logic_vector(x2_113 + to_signed(1,64))))) ) when others;

  x2_113 <= y_111;

  y_111 <= a1_54.Tup2_1_sel1_signed_1;

  a1_54 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_111\(127 downto 0)));

  -- index begin
  indexVec_111 : block
    signal vec_index_111 : integer range 0 to 64-1;
  begin
    vec_index_111 <= to_integer(resPtr_55)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_111\ <= currRes_55(vec_index_111);
  end block;
  -- index end

  currRes_55 <= \c$countConOut_app_arg_55\.Tup2_0_sel1_array_of_Maybe;

  resPtr_55 <= \c$countConOut_app_arg_55\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_112\ <= tagToEnum(\c$~<~Out_app_arg_113\);

  \c$~<~Out_app_arg_113\ <= to_signed(1,64) when x1_55 /= y_112 else to_signed(0,64);

  y_112 <= wild2_56;

  x1_55 <= wild2_55;

  -- index begin
  indexVec_112 : block
    signal vec_index_112 : integer range 0 to 64-1;
  begin
    vec_index_112 <= to_integer(to_signed(7,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_55 <= \c$app_arg\(vec_index_112);
  end block;
  -- index end

  \c$countConOut_app_arg_55\ <= ( Tup2_0_sel0_signed => x2_114 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_56\ ) when \c$~<~Out_case_scrut_114\ else
                                ( Tup2_0_sel0_signed => resPtr_56
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_56\ );

  clash_internal_cOut_56 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_56\
      , xs           => currRes_56
      , ds           => \c$~<~Out_app_arg_114\ );

  \c$~<~Out_app_arg_114\ <= ( Tup2_sel0_signed => x2_114 + to_signed(1,64)
                            , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_56)
                             & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_114\ else
                            \c$~<~Out_case_alt_55\;

  x2_114 <= resPtr_56;

  with (\c$~<~Out_case_scrut_113\(128 downto 128)) select
    \c$~<~Out_case_alt_55\ <= ( Tup2_sel0_signed => resPtr_56
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_57)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_56
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_57)
                               & std_logic_vector(x2_115 + to_signed(1,64))))) ) when others;

  x2_115 <= y_113;

  y_113 <= a1_55.Tup2_1_sel1_signed_1;

  a1_55 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_113\(127 downto 0)));

  -- index begin
  indexVec_113 : block
    signal vec_index_113 : integer range 0 to 64-1;
  begin
    vec_index_113 <= to_integer(resPtr_56)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_113\ <= currRes_56(vec_index_113);
  end block;
  -- index end

  currRes_56 <= \c$countConOut_app_arg_56\.Tup2_0_sel1_array_of_Maybe;

  resPtr_56 <= \c$countConOut_app_arg_56\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_114\ <= tagToEnum(\c$~<~Out_app_arg_115\);

  \c$~<~Out_app_arg_115\ <= to_signed(1,64) when x1_56 /= y_114 else to_signed(0,64);

  y_114 <= wild2_57;

  x1_56 <= wild2_56;

  -- index begin
  indexVec_114 : block
    signal vec_index_114 : integer range 0 to 64-1;
  begin
    vec_index_114 <= to_integer(to_signed(6,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_56 <= \c$app_arg\(vec_index_114);
  end block;
  -- index end

  \c$countConOut_app_arg_56\ <= ( Tup2_0_sel0_signed => x2_116 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_57\ ) when \c$~<~Out_case_scrut_116\ else
                                ( Tup2_0_sel0_signed => resPtr_57
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_57\ );

  clash_internal_cOut_57 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_57\
      , xs           => currRes_57
      , ds           => \c$~<~Out_app_arg_116\ );

  \c$~<~Out_app_arg_116\ <= ( Tup2_sel0_signed => x2_116 + to_signed(1,64)
                            , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_57)
                             & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_116\ else
                            \c$~<~Out_case_alt_56\;

  x2_116 <= resPtr_57;

  with (\c$~<~Out_case_scrut_115\(128 downto 128)) select
    \c$~<~Out_case_alt_56\ <= ( Tup2_sel0_signed => resPtr_57
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_58)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_57
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_58)
                               & std_logic_vector(x2_117 + to_signed(1,64))))) ) when others;

  x2_117 <= y_115;

  y_115 <= a1_56.Tup2_1_sel1_signed_1;

  a1_56 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_115\(127 downto 0)));

  -- index begin
  indexVec_115 : block
    signal vec_index_115 : integer range 0 to 64-1;
  begin
    vec_index_115 <= to_integer(resPtr_57)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_115\ <= currRes_57(vec_index_115);
  end block;
  -- index end

  currRes_57 <= \c$countConOut_app_arg_57\.Tup2_0_sel1_array_of_Maybe;

  resPtr_57 <= \c$countConOut_app_arg_57\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_116\ <= tagToEnum(\c$~<~Out_app_arg_117\);

  \c$~<~Out_app_arg_117\ <= to_signed(1,64) when x1_57 /= y_116 else to_signed(0,64);

  y_116 <= wild2_58;

  x1_57 <= wild2_57;

  -- index begin
  indexVec_116 : block
    signal vec_index_116 : integer range 0 to 64-1;
  begin
    vec_index_116 <= to_integer(to_signed(5,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_57 <= \c$app_arg\(vec_index_116);
  end block;
  -- index end

  \c$countConOut_app_arg_57\ <= ( Tup2_0_sel0_signed => x2_118 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_58\ ) when \c$~<~Out_case_scrut_118\ else
                                ( Tup2_0_sel0_signed => resPtr_58
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_58\ );

  clash_internal_cOut_58 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_58\
      , xs           => currRes_58
      , ds           => \c$~<~Out_app_arg_118\ );

  \c$~<~Out_app_arg_118\ <= ( Tup2_sel0_signed => x2_118 + to_signed(1,64)
                            , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_58)
                             & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_118\ else
                            \c$~<~Out_case_alt_57\;

  x2_118 <= resPtr_58;

  with (\c$~<~Out_case_scrut_117\(128 downto 128)) select
    \c$~<~Out_case_alt_57\ <= ( Tup2_sel0_signed => resPtr_58
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_59)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_58
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_59)
                               & std_logic_vector(x2_119 + to_signed(1,64))))) ) when others;

  x2_119 <= y_117;

  y_117 <= a1_57.Tup2_1_sel1_signed_1;

  a1_57 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_117\(127 downto 0)));

  -- index begin
  indexVec_117 : block
    signal vec_index_117 : integer range 0 to 64-1;
  begin
    vec_index_117 <= to_integer(resPtr_58)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_117\ <= currRes_58(vec_index_117);
  end block;
  -- index end

  currRes_58 <= \c$countConOut_app_arg_58\.Tup2_0_sel1_array_of_Maybe;

  resPtr_58 <= \c$countConOut_app_arg_58\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_118\ <= tagToEnum(\c$~<~Out_app_arg_119\);

  \c$~<~Out_app_arg_119\ <= to_signed(1,64) when x1_58 /= y_118 else to_signed(0,64);

  y_118 <= wild2_59;

  x1_58 <= wild2_58;

  -- index begin
  indexVec_118 : block
    signal vec_index_118 : integer range 0 to 64-1;
  begin
    vec_index_118 <= to_integer(to_signed(4,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_58 <= \c$app_arg\(vec_index_118);
  end block;
  -- index end

  \c$countConOut_app_arg_58\ <= ( Tup2_0_sel0_signed => x2_120 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_59\ ) when \c$~<~Out_case_scrut_120\ else
                                ( Tup2_0_sel0_signed => resPtr_59
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_59\ );

  clash_internal_cOut_59 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_59\
      , xs           => currRes_59
      , ds           => \c$~<~Out_app_arg_120\ );

  \c$~<~Out_app_arg_120\ <= ( Tup2_sel0_signed => x2_120 + to_signed(1,64)
                            , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_59)
                             & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_120\ else
                            \c$~<~Out_case_alt_58\;

  x2_120 <= resPtr_59;

  with (\c$~<~Out_case_scrut_119\(128 downto 128)) select
    \c$~<~Out_case_alt_58\ <= ( Tup2_sel0_signed => resPtr_59
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_60)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_59
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_60)
                               & std_logic_vector(x2_121 + to_signed(1,64))))) ) when others;

  x2_121 <= y_119;

  y_119 <= a1_58.Tup2_1_sel1_signed_1;

  a1_58 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_119\(127 downto 0)));

  -- index begin
  indexVec_119 : block
    signal vec_index_119 : integer range 0 to 64-1;
  begin
    vec_index_119 <= to_integer(resPtr_59)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_119\ <= currRes_59(vec_index_119);
  end block;
  -- index end

  currRes_59 <= \c$countConOut_app_arg_59\.Tup2_0_sel1_array_of_Maybe;

  resPtr_59 <= \c$countConOut_app_arg_59\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_120\ <= tagToEnum(\c$~<~Out_app_arg_121\);

  \c$~<~Out_app_arg_121\ <= to_signed(1,64) when x1_59 /= y_120 else to_signed(0,64);

  y_120 <= wild2_60;

  x1_59 <= wild2_59;

  -- index begin
  indexVec_120 : block
    signal vec_index_120 : integer range 0 to 64-1;
  begin
    vec_index_120 <= to_integer(to_signed(3,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_59 <= \c$app_arg\(vec_index_120);
  end block;
  -- index end

  \c$countConOut_app_arg_59\ <= ( Tup2_0_sel0_signed => x2_122 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_60\ ) when \c$~<~Out_case_scrut_122\ else
                                ( Tup2_0_sel0_signed => resPtr_60
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_60\ );

  clash_internal_cOut_60 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_60\
      , xs           => currRes_60
      , ds           => \c$~<~Out_app_arg_122\ );

  \c$~<~Out_app_arg_122\ <= ( Tup2_sel0_signed => x2_122 + to_signed(1,64)
                            , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_60)
                             & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_122\ else
                            \c$~<~Out_case_alt_59\;

  x2_122 <= resPtr_60;

  with (\c$~<~Out_case_scrut_121\(128 downto 128)) select
    \c$~<~Out_case_alt_59\ <= ( Tup2_sel0_signed => resPtr_60
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_61)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_60
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_61)
                               & std_logic_vector(x2_123 + to_signed(1,64))))) ) when others;

  x2_123 <= y_121;

  y_121 <= a1_59.Tup2_1_sel1_signed_1;

  a1_59 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_121\(127 downto 0)));

  -- index begin
  indexVec_121 : block
    signal vec_index_121 : integer range 0 to 64-1;
  begin
    vec_index_121 <= to_integer(resPtr_60)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_121\ <= currRes_60(vec_index_121);
  end block;
  -- index end

  currRes_60 <= \c$countConOut_app_arg_60\.Tup2_0_sel1_array_of_Maybe;

  resPtr_60 <= \c$countConOut_app_arg_60\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_122\ <= tagToEnum(\c$~<~Out_app_arg_123\);

  \c$~<~Out_app_arg_123\ <= to_signed(1,64) when x1_60 /= y_122 else to_signed(0,64);

  y_122 <= wild2_61;

  x1_60 <= wild2_60;

  -- index begin
  indexVec_122 : block
    signal vec_index_122 : integer range 0 to 64-1;
  begin
    vec_index_122 <= to_integer(to_signed(2,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_60 <= \c$app_arg\(vec_index_122);
  end block;
  -- index end

  \c$countConOut_app_arg_60\ <= ( Tup2_0_sel0_signed => x2_124 + to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_61\ ) when \c$~<~Out_case_scrut_124\ else
                                ( Tup2_0_sel0_signed => resPtr_61
                                , Tup2_0_sel1_array_of_Maybe => \c$~<~Out_61\ );

  clash_internal_cOut_61 : entity clash_internal
    port map
      ( \c$case_alt\ => \c$~<~Out_61\
      , xs           => currRes_61
      , ds           => \c$~<~Out_app_arg_124\ );

  \c$~<~Out_app_arg_124\ <= ( Tup2_sel0_signed => x2_124 + to_signed(1,64)
                            , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_61)
                             & std_logic_vector(to_signed(1,64))))) ) when \c$~<~Out_case_scrut_124\ else
                            \c$~<~Out_case_alt_60\;

  x2_124 <= resPtr_61;

  with (\c$~<~Out_case_scrut_123\(128 downto 128)) select
    \c$~<~Out_case_alt_60\ <= ( Tup2_sel0_signed => resPtr_61
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_62)
                               & std_logic_vector(to_signed(1,64))))) ) when "0",
                              ( Tup2_sel0_signed => resPtr_61
                              , Tup2_sel1_Maybe => std_logic_vector'("1" & ((std_logic_vector(wild2_62)
                               & std_logic_vector(x2_125 + to_signed(1,64))))) ) when others;

  x2_125 <= y_123;

  y_123 <= a1_60.Tup2_1_sel1_signed_1;

  a1_60 <= Main_topEntity_types.Tup2_1'(main_topentity_types.fromSLV(\c$~<~Out_case_scrut_123\(127 downto 0)));

  -- index begin
  indexVec_123 : block
    signal vec_index_123 : integer range 0 to 64-1;
  begin
    vec_index_123 <= to_integer(resPtr_61)
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    \c$~<~Out_case_scrut_123\ <= currRes_61(vec_index_123);
  end block;
  -- index end

  currRes_61 <= \c$countConOut_app_arg_62\.Tup2_0_sel1_array_of_Maybe;

  resPtr_61 <= \c$countConOut_app_arg_62\.Tup2_0_sel0_signed;

  \c$~<~Out_case_scrut_124\ <= tagToEnum(\c$~<~Out_app_arg_125\);

  \c$~<~Out_app_arg_125\ <= to_signed(1,64) when x1_61 /= y_124 else to_signed(0,64);

  y_124 <= wild2_62;

  x1_61 <= wild2_61;

  -- index begin
  indexVec_124 : block
    signal vec_index_124 : integer range 0 to 64-1;
  begin
    vec_index_124 <= to_integer(to_signed(1,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_61 <= \c$app_arg\(vec_index_124);
  end block;
  -- index end

  \c$countConOut_app_arg_61\ <= to_signed(1,64) when x1_62 /= to_signed(1,64) else to_signed(0,64);

  clash_internal_0_result_129 : entity clash_internal_0
    port map
      ( result                  => result_129
      , \c$countConOut_bindCsr\ => wild2_62 );

  \c$countConOut_case_scrut\ <= tagToEnum(\c$countConOut_app_arg_61\);

  \c$countConOut_app_arg_62\ <= ( Tup2_0_sel0_signed => to_signed(1,64)
                                , Tup2_0_sel1_array_of_Maybe => result_129 ) when \c$countConOut_case_scrut\ else
                                ( Tup2_0_sel0_signed => to_signed(0,64)
                                , Tup2_0_sel1_array_of_Maybe => Main_topEntity_types.array_of_Maybe'( std_logic_vector'("1" & ((std_logic_vector(to_signed(1,64))
                                                                                                     & std_logic_vector(to_signed(1,64)))))
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                                                                                    , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------") ) );

  -- index begin
  indexVec_125 : block
    signal vec_index_125 : integer range 0 to 64-1;
  begin
    vec_index_125 <= to_integer(to_signed(0,64))
    -- pragma translate_off
                 mod 64
    -- pragma translate_on
                 ;
    wild2_62 <= \c$app_arg\(vec_index_125);
  end block;
  -- index end

  x1_62 <= wild2_62;

  result <= result_128.Tup2_0_sel1_array_of_Maybe;

  result_0 <= result(0);

  result_1 <= result(1);

  result_2 <= result(2);

  result_3 <= result(3);

  result_4 <= result(4);

  result_5 <= result(5);

  result_6 <= result(6);

  result_7 <= result(7);

  result_8 <= result(8);

  result_9 <= result(9);

  result_10 <= result(10);

  result_11 <= result(11);

  result_12 <= result(12);

  result_13 <= result(13);

  result_14 <= result(14);

  result_15 <= result(15);

  result_16 <= result(16);

  result_17 <= result(17);

  result_18 <= result(18);

  result_19 <= result(19);

  result_20 <= result(20);

  result_21 <= result(21);

  result_22 <= result(22);

  result_23 <= result(23);

  result_24 <= result(24);

  result_25 <= result(25);

  result_26 <= result(26);

  result_27 <= result(27);

  result_28 <= result(28);

  result_29 <= result(29);

  result_30 <= result(30);

  result_31 <= result(31);

  result_32 <= result(32);

  result_33 <= result(33);

  result_34 <= result(34);

  result_35 <= result(35);

  result_36 <= result(36);

  result_37 <= result(37);

  result_38 <= result(38);

  result_39 <= result(39);

  result_40 <= result(40);

  result_41 <= result(41);

  result_42 <= result(42);

  result_43 <= result(43);

  result_44 <= result(44);

  result_45 <= result(45);

  result_46 <= result(46);

  result_47 <= result(47);

  result_48 <= result(48);

  result_49 <= result(49);

  result_50 <= result(50);

  result_51 <= result(51);

  result_52 <= result(52);

  result_53 <= result(53);

  result_54 <= result(54);

  result_55 <= result(55);

  result_56 <= result(56);

  result_57 <= result(57);

  result_58 <= result(58);

  result_59 <= result(59);

  result_60 <= result(60);

  result_61 <= result(61);

  result_62 <= result(62);

  result_63 <= result(63);


end;

