-- Automatically generated VHDL-93
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;
use std.textio.all;
use work.all;
use work.Main_topEntity_types.all;

entity matrixTraversalZigZag1 is
  port(\input\ : in Main_topEntity_types.array_of_array_of_8_signed_64(0 to 7);
       result  : out Main_topEntity_types.array_of_signed_64(0 to 63));
end;

architecture structural of matrixTraversalZigZag1 is
  signal \c$app_arg\    : signed(63 downto 0);
  signal \c$app_arg_0\  : signed(63 downto 0);
  signal \c$app_arg_1\  : signed(63 downto 0);
  signal \c$app_arg_2\  : signed(63 downto 0);
  signal \c$app_arg_3\  : signed(63 downto 0);
  signal \c$app_arg_4\  : signed(63 downto 0);
  signal \c$app_arg_5\  : signed(63 downto 0);
  signal \c$app_arg_6\  : signed(63 downto 0);
  signal \c$app_arg_7\  : signed(63 downto 0);
  signal \c$app_arg_8\  : signed(63 downto 0);
  signal \c$app_arg_9\  : signed(63 downto 0);
  signal \c$app_arg_10\ : signed(63 downto 0);
  signal \c$app_arg_11\ : signed(63 downto 0);
  signal \c$app_arg_12\ : signed(63 downto 0);
  signal \c$app_arg_13\ : signed(63 downto 0);
  signal \c$app_arg_14\ : signed(63 downto 0);
  signal \c$app_arg_15\ : signed(63 downto 0);
  signal \c$app_arg_16\ : signed(63 downto 0);
  signal \c$app_arg_17\ : signed(63 downto 0);
  signal \c$app_arg_18\ : signed(63 downto 0);
  signal \c$app_arg_19\ : signed(63 downto 0);
  signal \c$app_arg_20\ : signed(63 downto 0);
  signal \c$app_arg_21\ : signed(63 downto 0);
  signal \c$app_arg_22\ : signed(63 downto 0);
  signal \c$app_arg_23\ : signed(63 downto 0);
  signal \c$app_arg_24\ : signed(63 downto 0);
  signal \c$app_arg_25\ : signed(63 downto 0);
  signal \c$app_arg_26\ : signed(63 downto 0);
  signal \c$app_arg_27\ : signed(63 downto 0);
  signal \c$app_arg_28\ : Main_topEntity_types.array_of_signed_64(0 to 7);
  signal \c$app_arg_29\ : signed(63 downto 0);
  signal \c$app_arg_30\ : signed(63 downto 0);
  signal \c$app_arg_31\ : signed(63 downto 0);
  signal \c$app_arg_32\ : signed(63 downto 0);
  signal \c$app_arg_33\ : signed(63 downto 0);
  signal \c$app_arg_34\ : signed(63 downto 0);
  signal \c$app_arg_35\ : signed(63 downto 0);
  signal \c$app_arg_36\ : signed(63 downto 0);
  signal \c$app_arg_37\ : signed(63 downto 0);
  signal \c$app_arg_38\ : signed(63 downto 0);
  signal \c$app_arg_39\ : signed(63 downto 0);
  signal \c$app_arg_40\ : signed(63 downto 0);
  signal \c$app_arg_41\ : signed(63 downto 0);
  signal \c$app_arg_42\ : signed(63 downto 0);
  signal \c$app_arg_43\ : Main_topEntity_types.array_of_signed_64(0 to 7);
  signal \c$app_arg_44\ : signed(63 downto 0);
  signal \c$app_arg_45\ : Main_topEntity_types.array_of_signed_64(0 to 7);
  signal \c$app_arg_46\ : signed(63 downto 0);
  signal \c$app_arg_47\ : signed(63 downto 0);
  signal \c$app_arg_48\ : signed(63 downto 0);
  signal \c$app_arg_49\ : signed(63 downto 0);
  signal \c$app_arg_50\ : signed(63 downto 0);
  signal \c$app_arg_51\ : signed(63 downto 0);
  signal \c$app_arg_52\ : signed(63 downto 0);
  signal \c$app_arg_53\ : signed(63 downto 0);
  signal \c$app_arg_54\ : signed(63 downto 0);
  signal \c$app_arg_55\ : signed(63 downto 0);
  signal \c$app_arg_56\ : Main_topEntity_types.array_of_signed_64(0 to 7);
  signal \c$app_arg_57\ : signed(63 downto 0);
  signal \c$app_arg_58\ : Main_topEntity_types.array_of_signed_64(0 to 7);
  signal \c$app_arg_59\ : signed(63 downto 0);
  signal \c$app_arg_60\ : signed(63 downto 0);
  signal \c$app_arg_61\ : signed(63 downto 0);
  signal \c$app_arg_62\ : signed(63 downto 0);
  signal \c$app_arg_63\ : signed(63 downto 0);
  signal \c$app_arg_64\ : signed(63 downto 0);
  signal \c$app_arg_65\ : Main_topEntity_types.array_of_signed_64(0 to 7);
  signal \c$app_arg_66\ : signed(63 downto 0);
  signal \c$app_arg_67\ : Main_topEntity_types.array_of_signed_64(0 to 7);
  signal \c$app_arg_68\ : signed(63 downto 0);
  signal \c$app_arg_69\ : signed(63 downto 0);
  signal \c$app_arg_70\ : Main_topEntity_types.array_of_signed_64(0 to 7);

begin
  result <= Main_topEntity_types.array_of_signed_64'( \c$app_arg_69\
                                                    , \c$app_arg_68\
                                                    , \c$app_arg_66\
                                                    , \c$app_arg_64\
                                                    , \c$app_arg_63\
                                                    , \c$app_arg_62\
                                                    , \c$app_arg_61\
                                                    , \c$app_arg_60\
                                                    , \c$app_arg_59\
                                                    , \c$app_arg_57\
                                                    , \c$app_arg_55\
                                                    , \c$app_arg_54\
                                                    , \c$app_arg_53\
                                                    , \c$app_arg_52\
                                                    , \c$app_arg_51\
                                                    , \c$app_arg_50\
                                                    , \c$app_arg_49\
                                                    , \c$app_arg_48\
                                                    , \c$app_arg_47\
                                                    , \c$app_arg_46\
                                                    , \c$app_arg_44\
                                                    , \c$app_arg_42\
                                                    , \c$app_arg_41\
                                                    , \c$app_arg_40\
                                                    , \c$app_arg_39\
                                                    , \c$app_arg_38\
                                                    , \c$app_arg_37\
                                                    , \c$app_arg_36\
                                                    , \c$app_arg_35\
                                                    , \c$app_arg_34\
                                                    , \c$app_arg_33\
                                                    , \c$app_arg_32\
                                                    , \c$app_arg_31\
                                                    , \c$app_arg_30\
                                                    , \c$app_arg_29\
                                                    , \c$app_arg_27\
                                                    , \c$app_arg_26\
                                                    , \c$app_arg_25\
                                                    , \c$app_arg_24\
                                                    , \c$app_arg_23\
                                                    , \c$app_arg_22\
                                                    , \c$app_arg_21\
                                                    , \c$app_arg_20\
                                                    , \c$app_arg_19\
                                                    , \c$app_arg_18\
                                                    , \c$app_arg_17\
                                                    , \c$app_arg_16\
                                                    , \c$app_arg_15\
                                                    , \c$app_arg_14\
                                                    , \c$app_arg_13\
                                                    , \c$app_arg_12\
                                                    , \c$app_arg_11\
                                                    , \c$app_arg_10\
                                                    , \c$app_arg_9\
                                                    , \c$app_arg_8\
                                                    , \c$app_arg_7\
                                                    , \c$app_arg_6\
                                                    , \c$app_arg_5\
                                                    , \c$app_arg_4\
                                                    , \c$app_arg_3\
                                                    , \c$app_arg_2\
                                                    , \c$app_arg_1\
                                                    , \c$app_arg_0\
                                                    , \c$app_arg\ );

  -- index begin
  indexVec : block
    signal vec_index : integer range 0 to 8-1;
  begin
    vec_index <= to_integer(to_signed(7,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg\ <= \c$app_arg_28\(vec_index);
  end block;
  -- index end

  -- index begin
  indexVec_0 : block
    signal vec_index_0 : integer range 0 to 8-1;
  begin
    vec_index_0 <= to_integer(to_signed(6,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_0\ <= \c$app_arg_28\(vec_index_0);
  end block;
  -- index end

  -- index begin
  indexVec_1 : block
    signal vec_index_1 : integer range 0 to 8-1;
  begin
    vec_index_1 <= to_integer(to_signed(7,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_1\ <= \c$app_arg_43\(vec_index_1);
  end block;
  -- index end

  -- index begin
  indexVec_2 : block
    signal vec_index_2 : integer range 0 to 8-1;
  begin
    vec_index_2 <= to_integer(to_signed(7,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_2\ <= \c$app_arg_45\(vec_index_2);
  end block;
  -- index end

  -- index begin
  indexVec_3 : block
    signal vec_index_3 : integer range 0 to 8-1;
  begin
    vec_index_3 <= to_integer(to_signed(6,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_3\ <= \c$app_arg_43\(vec_index_3);
  end block;
  -- index end

  -- index begin
  indexVec_4 : block
    signal vec_index_4 : integer range 0 to 8-1;
  begin
    vec_index_4 <= to_integer(to_signed(5,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_4\ <= \c$app_arg_28\(vec_index_4);
  end block;
  -- index end

  -- index begin
  indexVec_5 : block
    signal vec_index_5 : integer range 0 to 8-1;
  begin
    vec_index_5 <= to_integer(to_signed(4,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_5\ <= \c$app_arg_28\(vec_index_5);
  end block;
  -- index end

  -- index begin
  indexVec_6 : block
    signal vec_index_6 : integer range 0 to 8-1;
  begin
    vec_index_6 <= to_integer(to_signed(5,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_6\ <= \c$app_arg_43\(vec_index_6);
  end block;
  -- index end

  -- index begin
  indexVec_7 : block
    signal vec_index_7 : integer range 0 to 8-1;
  begin
    vec_index_7 <= to_integer(to_signed(6,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_7\ <= \c$app_arg_45\(vec_index_7);
  end block;
  -- index end

  -- index begin
  indexVec_8 : block
    signal vec_index_8 : integer range 0 to 8-1;
  begin
    vec_index_8 <= to_integer(to_signed(7,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_8\ <= \c$app_arg_56\(vec_index_8);
  end block;
  -- index end

  -- index begin
  indexVec_9 : block
    signal vec_index_9 : integer range 0 to 8-1;
  begin
    vec_index_9 <= to_integer(to_signed(7,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_9\ <= \c$app_arg_58\(vec_index_9);
  end block;
  -- index end

  -- index begin
  indexVec_10 : block
    signal vec_index_10 : integer range 0 to 8-1;
  begin
    vec_index_10 <= to_integer(to_signed(6,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_10\ <= \c$app_arg_56\(vec_index_10);
  end block;
  -- index end

  -- index begin
  indexVec_11 : block
    signal vec_index_11 : integer range 0 to 8-1;
  begin
    vec_index_11 <= to_integer(to_signed(5,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_11\ <= \c$app_arg_45\(vec_index_11);
  end block;
  -- index end

  -- index begin
  indexVec_12 : block
    signal vec_index_12 : integer range 0 to 8-1;
  begin
    vec_index_12 <= to_integer(to_signed(4,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_12\ <= \c$app_arg_43\(vec_index_12);
  end block;
  -- index end

  -- index begin
  indexVec_13 : block
    signal vec_index_13 : integer range 0 to 8-1;
  begin
    vec_index_13 <= to_integer(to_signed(3,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_13\ <= \c$app_arg_28\(vec_index_13);
  end block;
  -- index end

  -- index begin
  indexVec_14 : block
    signal vec_index_14 : integer range 0 to 8-1;
  begin
    vec_index_14 <= to_integer(to_signed(2,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_14\ <= \c$app_arg_28\(vec_index_14);
  end block;
  -- index end

  -- index begin
  indexVec_15 : block
    signal vec_index_15 : integer range 0 to 8-1;
  begin
    vec_index_15 <= to_integer(to_signed(3,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_15\ <= \c$app_arg_43\(vec_index_15);
  end block;
  -- index end

  -- index begin
  indexVec_16 : block
    signal vec_index_16 : integer range 0 to 8-1;
  begin
    vec_index_16 <= to_integer(to_signed(4,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_16\ <= \c$app_arg_45\(vec_index_16);
  end block;
  -- index end

  -- index begin
  indexVec_17 : block
    signal vec_index_17 : integer range 0 to 8-1;
  begin
    vec_index_17 <= to_integer(to_signed(5,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_17\ <= \c$app_arg_56\(vec_index_17);
  end block;
  -- index end

  -- index begin
  indexVec_18 : block
    signal vec_index_18 : integer range 0 to 8-1;
  begin
    vec_index_18 <= to_integer(to_signed(6,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_18\ <= \c$app_arg_58\(vec_index_18);
  end block;
  -- index end

  -- index begin
  indexVec_19 : block
    signal vec_index_19 : integer range 0 to 8-1;
  begin
    vec_index_19 <= to_integer(to_signed(7,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_19\ <= \c$app_arg_65\(vec_index_19);
  end block;
  -- index end

  -- index begin
  indexVec_20 : block
    signal vec_index_20 : integer range 0 to 8-1;
  begin
    vec_index_20 <= to_integer(to_signed(7,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_20\ <= \c$app_arg_67\(vec_index_20);
  end block;
  -- index end

  -- index begin
  indexVec_21 : block
    signal vec_index_21 : integer range 0 to 8-1;
  begin
    vec_index_21 <= to_integer(to_signed(6,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_21\ <= \c$app_arg_65\(vec_index_21);
  end block;
  -- index end

  -- index begin
  indexVec_22 : block
    signal vec_index_22 : integer range 0 to 8-1;
  begin
    vec_index_22 <= to_integer(to_signed(5,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_22\ <= \c$app_arg_58\(vec_index_22);
  end block;
  -- index end

  -- index begin
  indexVec_23 : block
    signal vec_index_23 : integer range 0 to 8-1;
  begin
    vec_index_23 <= to_integer(to_signed(4,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_23\ <= \c$app_arg_56\(vec_index_23);
  end block;
  -- index end

  -- index begin
  indexVec_24 : block
    signal vec_index_24 : integer range 0 to 8-1;
  begin
    vec_index_24 <= to_integer(to_signed(3,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_24\ <= \c$app_arg_45\(vec_index_24);
  end block;
  -- index end

  -- index begin
  indexVec_25 : block
    signal vec_index_25 : integer range 0 to 8-1;
  begin
    vec_index_25 <= to_integer(to_signed(2,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_25\ <= \c$app_arg_43\(vec_index_25);
  end block;
  -- index end

  -- index begin
  indexVec_26 : block
    signal vec_index_26 : integer range 0 to 8-1;
  begin
    vec_index_26 <= to_integer(to_signed(1,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_26\ <= \c$app_arg_28\(vec_index_26);
  end block;
  -- index end

  -- index begin
  indexVec_27 : block
    signal vec_index_27 : integer range 0 to 8-1;
  begin
    vec_index_27 <= to_integer(to_signed(0,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_27\ <= \c$app_arg_28\(vec_index_27);
  end block;
  -- index end

  -- index begin
  indexVec_28 : block
    signal vec_index_28 : integer range 0 to 8-1;
  begin
    vec_index_28 <= to_integer(to_signed(7,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_28\ <= \input\(vec_index_28);
  end block;
  -- index end

  -- index begin
  indexVec_29 : block
    signal vec_index_29 : integer range 0 to 8-1;
  begin
    vec_index_29 <= to_integer(to_signed(1,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_29\ <= \c$app_arg_43\(vec_index_29);
  end block;
  -- index end

  -- index begin
  indexVec_30 : block
    signal vec_index_30 : integer range 0 to 8-1;
  begin
    vec_index_30 <= to_integer(to_signed(2,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_30\ <= \c$app_arg_45\(vec_index_30);
  end block;
  -- index end

  -- index begin
  indexVec_31 : block
    signal vec_index_31 : integer range 0 to 8-1;
  begin
    vec_index_31 <= to_integer(to_signed(3,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_31\ <= \c$app_arg_56\(vec_index_31);
  end block;
  -- index end

  -- index begin
  indexVec_32 : block
    signal vec_index_32 : integer range 0 to 8-1;
  begin
    vec_index_32 <= to_integer(to_signed(4,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_32\ <= \c$app_arg_58\(vec_index_32);
  end block;
  -- index end

  -- index begin
  indexVec_33 : block
    signal vec_index_33 : integer range 0 to 8-1;
  begin
    vec_index_33 <= to_integer(to_signed(5,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_33\ <= \c$app_arg_65\(vec_index_33);
  end block;
  -- index end

  -- index begin
  indexVec_34 : block
    signal vec_index_34 : integer range 0 to 8-1;
  begin
    vec_index_34 <= to_integer(to_signed(6,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_34\ <= \c$app_arg_67\(vec_index_34);
  end block;
  -- index end

  -- index begin
  indexVec_35 : block
    signal vec_index_35 : integer range 0 to 8-1;
  begin
    vec_index_35 <= to_integer(to_signed(7,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_35\ <= \c$app_arg_70\(vec_index_35);
  end block;
  -- index end

  -- index begin
  indexVec_36 : block
    signal vec_index_36 : integer range 0 to 8-1;
  begin
    vec_index_36 <= to_integer(to_signed(6,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_36\ <= \c$app_arg_70\(vec_index_36);
  end block;
  -- index end

  -- index begin
  indexVec_37 : block
    signal vec_index_37 : integer range 0 to 8-1;
  begin
    vec_index_37 <= to_integer(to_signed(5,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_37\ <= \c$app_arg_67\(vec_index_37);
  end block;
  -- index end

  -- index begin
  indexVec_38 : block
    signal vec_index_38 : integer range 0 to 8-1;
  begin
    vec_index_38 <= to_integer(to_signed(4,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_38\ <= \c$app_arg_65\(vec_index_38);
  end block;
  -- index end

  -- index begin
  indexVec_39 : block
    signal vec_index_39 : integer range 0 to 8-1;
  begin
    vec_index_39 <= to_integer(to_signed(3,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_39\ <= \c$app_arg_58\(vec_index_39);
  end block;
  -- index end

  -- index begin
  indexVec_40 : block
    signal vec_index_40 : integer range 0 to 8-1;
  begin
    vec_index_40 <= to_integer(to_signed(2,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_40\ <= \c$app_arg_56\(vec_index_40);
  end block;
  -- index end

  -- index begin
  indexVec_41 : block
    signal vec_index_41 : integer range 0 to 8-1;
  begin
    vec_index_41 <= to_integer(to_signed(1,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_41\ <= \c$app_arg_45\(vec_index_41);
  end block;
  -- index end

  -- index begin
  indexVec_42 : block
    signal vec_index_42 : integer range 0 to 8-1;
  begin
    vec_index_42 <= to_integer(to_signed(0,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_42\ <= \c$app_arg_43\(vec_index_42);
  end block;
  -- index end

  -- index begin
  indexVec_43 : block
    signal vec_index_43 : integer range 0 to 8-1;
  begin
    vec_index_43 <= to_integer(to_signed(6,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_43\ <= \input\(vec_index_43);
  end block;
  -- index end

  -- index begin
  indexVec_44 : block
    signal vec_index_44 : integer range 0 to 8-1;
  begin
    vec_index_44 <= to_integer(to_signed(0,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_44\ <= \c$app_arg_45\(vec_index_44);
  end block;
  -- index end

  -- index begin
  indexVec_45 : block
    signal vec_index_45 : integer range 0 to 8-1;
  begin
    vec_index_45 <= to_integer(to_signed(5,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_45\ <= \input\(vec_index_45);
  end block;
  -- index end

  -- index begin
  indexVec_46 : block
    signal vec_index_46 : integer range 0 to 8-1;
  begin
    vec_index_46 <= to_integer(to_signed(1,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_46\ <= \c$app_arg_56\(vec_index_46);
  end block;
  -- index end

  -- index begin
  indexVec_47 : block
    signal vec_index_47 : integer range 0 to 8-1;
  begin
    vec_index_47 <= to_integer(to_signed(2,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_47\ <= \c$app_arg_58\(vec_index_47);
  end block;
  -- index end

  -- index begin
  indexVec_48 : block
    signal vec_index_48 : integer range 0 to 8-1;
  begin
    vec_index_48 <= to_integer(to_signed(3,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_48\ <= \c$app_arg_65\(vec_index_48);
  end block;
  -- index end

  -- index begin
  indexVec_49 : block
    signal vec_index_49 : integer range 0 to 8-1;
  begin
    vec_index_49 <= to_integer(to_signed(4,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_49\ <= \c$app_arg_67\(vec_index_49);
  end block;
  -- index end

  -- index begin
  indexVec_50 : block
    signal vec_index_50 : integer range 0 to 8-1;
  begin
    vec_index_50 <= to_integer(to_signed(5,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_50\ <= \c$app_arg_70\(vec_index_50);
  end block;
  -- index end

  -- index begin
  indexVec_51 : block
    signal vec_index_51 : integer range 0 to 8-1;
  begin
    vec_index_51 <= to_integer(to_signed(4,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_51\ <= \c$app_arg_70\(vec_index_51);
  end block;
  -- index end

  -- index begin
  indexVec_52 : block
    signal vec_index_52 : integer range 0 to 8-1;
  begin
    vec_index_52 <= to_integer(to_signed(3,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_52\ <= \c$app_arg_67\(vec_index_52);
  end block;
  -- index end

  -- index begin
  indexVec_53 : block
    signal vec_index_53 : integer range 0 to 8-1;
  begin
    vec_index_53 <= to_integer(to_signed(2,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_53\ <= \c$app_arg_65\(vec_index_53);
  end block;
  -- index end

  -- index begin
  indexVec_54 : block
    signal vec_index_54 : integer range 0 to 8-1;
  begin
    vec_index_54 <= to_integer(to_signed(1,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_54\ <= \c$app_arg_58\(vec_index_54);
  end block;
  -- index end

  -- index begin
  indexVec_55 : block
    signal vec_index_55 : integer range 0 to 8-1;
  begin
    vec_index_55 <= to_integer(to_signed(0,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_55\ <= \c$app_arg_56\(vec_index_55);
  end block;
  -- index end

  -- index begin
  indexVec_56 : block
    signal vec_index_56 : integer range 0 to 8-1;
  begin
    vec_index_56 <= to_integer(to_signed(4,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_56\ <= \input\(vec_index_56);
  end block;
  -- index end

  -- index begin
  indexVec_57 : block
    signal vec_index_57 : integer range 0 to 8-1;
  begin
    vec_index_57 <= to_integer(to_signed(0,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_57\ <= \c$app_arg_58\(vec_index_57);
  end block;
  -- index end

  -- index begin
  indexVec_58 : block
    signal vec_index_58 : integer range 0 to 8-1;
  begin
    vec_index_58 <= to_integer(to_signed(3,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_58\ <= \input\(vec_index_58);
  end block;
  -- index end

  -- index begin
  indexVec_59 : block
    signal vec_index_59 : integer range 0 to 8-1;
  begin
    vec_index_59 <= to_integer(to_signed(1,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_59\ <= \c$app_arg_65\(vec_index_59);
  end block;
  -- index end

  -- index begin
  indexVec_60 : block
    signal vec_index_60 : integer range 0 to 8-1;
  begin
    vec_index_60 <= to_integer(to_signed(2,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_60\ <= \c$app_arg_67\(vec_index_60);
  end block;
  -- index end

  -- index begin
  indexVec_61 : block
    signal vec_index_61 : integer range 0 to 8-1;
  begin
    vec_index_61 <= to_integer(to_signed(3,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_61\ <= \c$app_arg_70\(vec_index_61);
  end block;
  -- index end

  -- index begin
  indexVec_62 : block
    signal vec_index_62 : integer range 0 to 8-1;
  begin
    vec_index_62 <= to_integer(to_signed(2,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_62\ <= \c$app_arg_70\(vec_index_62);
  end block;
  -- index end

  -- index begin
  indexVec_63 : block
    signal vec_index_63 : integer range 0 to 8-1;
  begin
    vec_index_63 <= to_integer(to_signed(1,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_63\ <= \c$app_arg_67\(vec_index_63);
  end block;
  -- index end

  -- index begin
  indexVec_64 : block
    signal vec_index_64 : integer range 0 to 8-1;
  begin
    vec_index_64 <= to_integer(to_signed(0,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_64\ <= \c$app_arg_65\(vec_index_64);
  end block;
  -- index end

  -- index begin
  indexVec_65 : block
    signal vec_index_65 : integer range 0 to 8-1;
  begin
    vec_index_65 <= to_integer(to_signed(2,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_65\ <= \input\(vec_index_65);
  end block;
  -- index end

  -- index begin
  indexVec_66 : block
    signal vec_index_66 : integer range 0 to 8-1;
  begin
    vec_index_66 <= to_integer(to_signed(0,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_66\ <= \c$app_arg_67\(vec_index_66);
  end block;
  -- index end

  -- index begin
  indexVec_67 : block
    signal vec_index_67 : integer range 0 to 8-1;
  begin
    vec_index_67 <= to_integer(to_signed(1,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_67\ <= \input\(vec_index_67);
  end block;
  -- index end

  -- index begin
  indexVec_68 : block
    signal vec_index_68 : integer range 0 to 8-1;
  begin
    vec_index_68 <= to_integer(to_signed(1,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_68\ <= \c$app_arg_70\(vec_index_68);
  end block;
  -- index end

  -- index begin
  indexVec_69 : block
    signal vec_index_69 : integer range 0 to 8-1;
  begin
    vec_index_69 <= to_integer(to_signed(0,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_69\ <= \c$app_arg_70\(vec_index_69);
  end block;
  -- index end

  -- index begin
  indexVec_70 : block
    signal vec_index_70 : integer range 0 to 8-1;
  begin
    vec_index_70 <= to_integer(to_signed(0,64))
    -- pragma translate_off
                 mod 8
    -- pragma translate_on
                 ;
    \c$app_arg_70\ <= \input\(vec_index_70);
  end block;
  -- index end


end;

