-- Automatically generated VHDL-93
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;
use std.textio.all;
use work.all;
use work.Main_topEntity_types.all;

entity clash_internal_0 is
  port(\c$countConOut_bindCsr\ : in signed(63 downto 0);
       result                  : out Main_topEntity_types.array_of_Maybe(0 to 63));
end;

architecture structural of clash_internal_0 is
  signal \result__dc_arg_res\ : Main_topEntity_types.array_of_Maybe(0 to 62);

begin
  -- replace begin
  replaceVec : block
    signal vec_index : integer range 0 to 63-1;
  begin
    vec_index <= to_integer(to_signed(0,64))
    -- pragma translate_off
                 mod 63
    -- pragma translate_on
                 ;

    process(vec_index,\c$countConOut_bindCsr\)
      variable ivec : Main_topEntity_types.array_of_Maybe(0 to 62);
    begin
      ivec := Main_topEntity_types.array_of_Maybe'( std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")
                                      , std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------") );
      ivec(vec_index) := std_logic_vector'("1" & ((std_logic_vector(\c$countConOut_bindCsr\)
   & std_logic_vector(to_signed(1,64)))));
      \result__dc_arg_res\ <= ivec;
    end process;
  end block;
  -- replace end

  result <= Main_topEntity_types.array_of_Maybe'(Main_topEntity_types.Maybe'(std_logic_vector'("0" & "--------------------------------------------------------------------------------------------------------------------------------")) & \result__dc_arg_res\);


end;

